module tt_um_julke_gussinatorn2
  (input  [7:0] ui_in,
   input  [7:0] uio_in,
   input  ena,
   input  clk,
   input  rst_n,
   output [7:0] uo_out,
   output [7:0] uio_out,
   output [7:0] uio_oe);
  reg [255:0] rom_mrse;
  reg [1:0] ascell_mrse;
  reg [1:0] cell_mrse;
  reg [5:0] ui_in_old;
  reg [5:0] ui_in_sync;
  reg [7:0] sr_mrse;
  reg [2:0] i_sr_mrse;
  reg flush_sr_mrse;
  reg [4:0] i_rom_mrse;
  reg [13:0] time_mrse;
  reg [2:0] state_mrse;
  localparam [7:0] n14_o = 8'b00000000;
  localparam [7:0] n15_o = 8'b00000000;
  wire [5:0] n16_o;
  wire [5:0] n17_o;
  wire [5:0] n18_o;
  wire n21_o;
  wire n22_o;
  wire n23_o;
  wire n24_o;
  wire n25_o;
  wire [1:0] n26_o;
  wire [1:0] n28_o;
  wire [5:0] n33_o;
  wire n35_o;
  wire n36_o;
  wire n38_o;
  wire n40_o;
  wire [31:0] n43_o;
  wire [31:0] n45_o;
  wire [4:0] n46_o;
  wire n47_o;
  wire n48_o;
  wire n49_o;
  wire n50_o;
  wire [5:0] n51_o;
  wire [7:0] n52_o;
  wire [2:0] n54_o;
  wire [7:0] n55_o;
  wire [2:0] n56_o;
  wire [255:0] n57_o;
  wire [7:0] n59_o;
  wire [2:0] n61_o;
  wire n63_o;
  wire [4:0] n64_o;
  wire n65_o;
  wire [7:0] n66_o;
  wire [2:0] n67_o;
  wire n69_o;
  wire n70_o;
  wire n71_o;
  wire n72_o;
  wire [2:0] n74_o;
  wire [4:0] n76_o;
  wire [2:0] n78_o;
  wire [2:0] n80_o;
  wire [4:0] n82_o;
  wire [2:0] n84_o;
  wire [2:0] n86_o;
  wire [4:0] n88_o;
  wire [2:0] n90_o;
  wire n92_o;
  wire [31:0] n93_o;
  wire n95_o;
  wire [2:0] n97_o;
  wire [4:0] n99_o;
  wire [2:0] n102_o;
  wire n104_o;
  wire [31:0] n105_o;
  wire [31:0] n107_o;
  wire [4:0] n108_o;
  wire [2:0] n110_o;
  wire [4:0] n111_o;
  wire [1:0] n114_o;
  wire n116_o;
  wire [1:0] n117_o;
  wire n119_o;
  wire [1:0] n120_o;
  wire n122_o;
  wire [1:0] n123_o;
  wire n125_o;
  wire [3:0] n126_o;
  reg [1:0] n127_o;
  wire n129_o;
  wire [31:0] n130_o;
  wire n132_o;
  wire [31:0] n133_o;
  wire [31:0] n135_o;
  wire [13:0] n136_o;
  wire [31:0] n138_o;
  wire n140_o;
  wire [31:0] n142_o;
  wire [31:0] n144_o;
  wire [13:0] n145_o;
  wire [2:0] n147_o;
  wire n148_o;
  wire n149_o;
  wire [2:0] n150_o;
  wire [13:0] n151_o;
  wire [2:0] n153_o;
  wire n154_o;
  wire [2:0] n155_o;
  wire [13:0] n156_o;
  wire [2:0] n157_o;
  wire n159_o;
  wire n163_o;
  wire [2:0] n165_o;
  wire [2:0] n166_o;
  wire n168_o;
  wire n172_o;
  wire [2:0] n174_o;
  wire [2:0] n175_o;
  wire n177_o;
  wire n179_o;
  wire n181_o;
  wire [3:0] n182_o;
  reg [7:0] n183_o;
  reg [2:0] n184_o;
  reg [13:0] n187_o;
  reg [2:0] n192_o;
  wire n194_o;
  wire [31:0] n195_o;
  wire n197_o;
  wire n200_o;
  wire [7:0] n202_o;
  wire [31:0] n204_o;
  wire [31:0] n206_o;
  wire [4:0] n207_o;
  wire [255:0] n210_o;
  wire [7:0] n211_o;
  wire [4:0] n212_o;
  wire n213_o;
  wire [7:0] n214_o;
  wire [4:0] n216_o;
  wire [2:0] n218_o;
  wire n220_o;
  wire [31:0] n221_o;
  wire n223_o;
  wire n226_o;
  wire [7:0] n228_o;
  wire [31:0] n230_o;
  wire [31:0] n232_o;
  wire [4:0] n233_o;
  wire [255:0] n236_o;
  wire [7:0] n237_o;
  wire [4:0] n238_o;
  wire n239_o;
  wire [7:0] n240_o;
  wire [4:0] n242_o;
  wire [2:0] n244_o;
  wire n245_o;
  wire n246_o;
  wire [4:0] n247_o;
  wire [2:0] n248_o;
  wire [255:0] n249_o;
  wire [7:0] n250_o;
  wire [4:0] n251_o;
  wire [2:0] n252_o;
  wire [255:0] n253_o;
  wire [7:0] n254_o;
  wire [2:0] n255_o;
  wire [4:0] n256_o;
  wire [13:0] n257_o;
  wire [2:0] n258_o;
  wire n259_o;
  wire n260_o;
  wire [255:0] n261_o;
  wire [7:0] n262_o;
  wire [2:0] n263_o;
  wire [4:0] n264_o;
  wire [13:0] n265_o;
  wire [2:0] n266_o;
  wire n267_o;
  wire n268_o;
  wire [255:0] n269_o;
  wire [7:0] n271_o;
  wire [2:0] n272_o;
  wire [4:0] n273_o;
  wire [13:0] n274_o;
  wire [2:0] n275_o;
  wire [6:0] n290_o;
  wire [6:0] n291_o;
  reg [255:0] n305_q;
  wire n306_o;
  wire n307_o;
  wire [1:0] n308_o;
  reg [1:0] n309_q;
  wire n310_o;
  wire [5:0] n311_o;
  reg [5:0] n312_q;
  wire n313_o;
  wire [7:0] n314_o;
  reg [7:0] n315_q;
  reg [2:0] n316_q;
  wire n317_o;
  wire n318_o;
  wire n319_o;
  reg n320_q;
  reg [4:0] n321_q;
  wire n322_o;
  wire [13:0] n323_o;
  reg [13:0] n324_q;
  wire n325_o;
  wire [2:0] n326_o;
  reg [2:0] n327_q;
  reg n328_q;
  wire [7:0] n329_o;
  wire n330_o;
  wire n331_o;
  wire n332_o;
  wire n333_o;
  wire n334_o;
  wire n335_o;
  wire n336_o;
  wire n337_o;
  wire n338_o;
  wire n339_o;
  wire n340_o;
  wire n341_o;
  wire n342_o;
  wire n343_o;
  wire n344_o;
  wire n345_o;
  wire n346_o;
  wire n347_o;
  wire n348_o;
  wire n349_o;
  wire n350_o;
  wire n351_o;
  wire n352_o;
  wire n353_o;
  wire n354_o;
  wire n355_o;
  wire n356_o;
  wire n357_o;
  wire n358_o;
  wire n359_o;
  wire n360_o;
  wire n361_o;
  wire n362_o;
  wire n363_o;
  wire n364_o;
  wire n365_o;
  wire n366_o;
  wire n367_o;
  wire n368_o;
  wire n369_o;
  wire n370_o;
  wire n371_o;
  wire n372_o;
  wire n373_o;
  wire n374_o;
  wire n375_o;
  wire n376_o;
  wire n377_o;
  wire n378_o;
  wire n379_o;
  wire n380_o;
  wire n381_o;
  wire n382_o;
  wire n383_o;
  wire n384_o;
  wire n385_o;
  wire n386_o;
  wire n387_o;
  wire n388_o;
  wire n389_o;
  wire n390_o;
  wire n391_o;
  wire n392_o;
  wire n393_o;
  wire n394_o;
  wire n395_o;
  wire n396_o;
  wire n397_o;
  wire n398_o;
  wire n399_o;
  wire [7:0] n400_o;
  wire [7:0] n401_o;
  wire [7:0] n402_o;
  wire [7:0] n403_o;
  wire [7:0] n404_o;
  wire [7:0] n405_o;
  wire [7:0] n406_o;
  wire [7:0] n407_o;
  wire [7:0] n408_o;
  wire [7:0] n409_o;
  wire [7:0] n410_o;
  wire [7:0] n411_o;
  wire [7:0] n412_o;
  wire [7:0] n413_o;
  wire [7:0] n414_o;
  wire [7:0] n415_o;
  wire [7:0] n416_o;
  wire [7:0] n417_o;
  wire [7:0] n418_o;
  wire [7:0] n419_o;
  wire [7:0] n420_o;
  wire [7:0] n421_o;
  wire [7:0] n422_o;
  wire [7:0] n423_o;
  wire [7:0] n424_o;
  wire [7:0] n425_o;
  wire [7:0] n426_o;
  wire [7:0] n427_o;
  wire [7:0] n428_o;
  wire [7:0] n429_o;
  wire [7:0] n430_o;
  wire [7:0] n431_o;
  wire [7:0] n432_o;
  wire [7:0] n433_o;
  wire [7:0] n434_o;
  wire [7:0] n435_o;
  wire [7:0] n436_o;
  wire [7:0] n437_o;
  wire [7:0] n438_o;
  wire [7:0] n439_o;
  wire [7:0] n440_o;
  wire [7:0] n441_o;
  wire [7:0] n442_o;
  wire [7:0] n443_o;
  wire [7:0] n444_o;
  wire [7:0] n445_o;
  wire [7:0] n446_o;
  wire [7:0] n447_o;
  wire [7:0] n448_o;
  wire [7:0] n449_o;
  wire [7:0] n450_o;
  wire [7:0] n451_o;
  wire [7:0] n452_o;
  wire [7:0] n453_o;
  wire [7:0] n454_o;
  wire [7:0] n455_o;
  wire [7:0] n456_o;
  wire [7:0] n457_o;
  wire [7:0] n458_o;
  wire [7:0] n459_o;
  wire [7:0] n460_o;
  wire [7:0] n461_o;
  wire [7:0] n462_o;
  wire [7:0] n463_o;
  wire [255:0] n464_o;
  wire [7:0] n465_o;
  wire [7:0] n466_o;
  wire [7:0] n467_o;
  wire [7:0] n468_o;
  wire [7:0] n469_o;
  wire [7:0] n470_o;
  wire [7:0] n471_o;
  wire [7:0] n472_o;
  wire [7:0] n473_o;
  wire [7:0] n474_o;
  wire [7:0] n475_o;
  wire [7:0] n476_o;
  wire [7:0] n477_o;
  wire [7:0] n478_o;
  wire [7:0] n479_o;
  wire [7:0] n480_o;
  wire [7:0] n481_o;
  wire [7:0] n482_o;
  wire [7:0] n483_o;
  wire [7:0] n484_o;
  wire [7:0] n485_o;
  wire [7:0] n486_o;
  wire [7:0] n487_o;
  wire [7:0] n488_o;
  wire [7:0] n489_o;
  wire [7:0] n490_o;
  wire [7:0] n491_o;
  wire [7:0] n492_o;
  wire [7:0] n493_o;
  wire [7:0] n494_o;
  wire [7:0] n495_o;
  wire [7:0] n496_o;
  wire [1:0] n497_o;
  reg [7:0] n498_o;
  wire [1:0] n499_o;
  reg [7:0] n500_o;
  wire [1:0] n501_o;
  reg [7:0] n502_o;
  wire [1:0] n503_o;
  reg [7:0] n504_o;
  wire [1:0] n505_o;
  reg [7:0] n506_o;
  wire [1:0] n507_o;
  reg [7:0] n508_o;
  wire [1:0] n509_o;
  reg [7:0] n510_o;
  wire [1:0] n511_o;
  reg [7:0] n512_o;
  wire [1:0] n513_o;
  reg [7:0] n514_o;
  wire [1:0] n515_o;
  reg [7:0] n516_o;
  wire n517_o;
  wire [7:0] n518_o;
  wire [7:0] n519_o;
  wire [7:0] n520_o;
  wire [7:0] n521_o;
  wire [7:0] n522_o;
  wire [7:0] n523_o;
  wire [7:0] n524_o;
  wire [7:0] n525_o;
  wire [7:0] n526_o;
  wire [7:0] n527_o;
  wire [7:0] n528_o;
  wire [7:0] n529_o;
  wire [7:0] n530_o;
  wire [7:0] n531_o;
  wire [7:0] n532_o;
  wire [7:0] n533_o;
  wire [7:0] n534_o;
  wire [7:0] n535_o;
  wire [7:0] n536_o;
  wire [7:0] n537_o;
  wire [7:0] n538_o;
  wire [7:0] n539_o;
  wire [7:0] n540_o;
  wire [7:0] n541_o;
  wire [7:0] n542_o;
  wire [7:0] n543_o;
  wire [7:0] n544_o;
  wire [7:0] n545_o;
  wire [7:0] n546_o;
  wire [7:0] n547_o;
  wire [7:0] n548_o;
  wire [7:0] n549_o;
  wire [7:0] n550_o;
  wire [1:0] n551_o;
  reg [7:0] n552_o;
  wire [1:0] n553_o;
  reg [7:0] n554_o;
  wire [1:0] n555_o;
  reg [7:0] n556_o;
  wire [1:0] n557_o;
  reg [7:0] n558_o;
  wire [1:0] n559_o;
  reg [7:0] n560_o;
  wire [1:0] n561_o;
  reg [7:0] n562_o;
  wire [1:0] n563_o;
  reg [7:0] n564_o;
  wire [1:0] n565_o;
  reg [7:0] n566_o;
  wire [1:0] n567_o;
  reg [7:0] n568_o;
  wire [1:0] n569_o;
  reg [7:0] n570_o;
  wire n571_o;
  wire [7:0] n572_o;
  wire [7:0] n573_o;
  wire [7:0] n574_o;
  wire [7:0] n575_o;
  wire [7:0] n576_o;
  wire [7:0] n577_o;
  wire [7:0] n578_o;
  wire [7:0] n579_o;
  wire [7:0] n580_o;
  wire [7:0] n581_o;
  wire [7:0] n582_o;
  wire [7:0] n583_o;
  wire [7:0] n584_o;
  wire [7:0] n585_o;
  wire [7:0] n586_o;
  wire [7:0] n587_o;
  wire [7:0] n588_o;
  wire [7:0] n589_o;
  wire [7:0] n590_o;
  wire [7:0] n591_o;
  wire [7:0] n592_o;
  wire [7:0] n593_o;
  wire [7:0] n594_o;
  wire [7:0] n595_o;
  wire [7:0] n596_o;
  wire [7:0] n597_o;
  wire [7:0] n598_o;
  wire [7:0] n599_o;
  wire [7:0] n600_o;
  wire [7:0] n601_o;
  wire [7:0] n602_o;
  wire [7:0] n603_o;
  wire [7:0] n604_o;
  wire [1:0] n605_o;
  reg [7:0] n606_o;
  wire [1:0] n607_o;
  reg [7:0] n608_o;
  wire [1:0] n609_o;
  reg [7:0] n610_o;
  wire [1:0] n611_o;
  reg [7:0] n612_o;
  wire [1:0] n613_o;
  reg [7:0] n614_o;
  wire [1:0] n615_o;
  reg [7:0] n616_o;
  wire [1:0] n617_o;
  reg [7:0] n618_o;
  wire [1:0] n619_o;
  reg [7:0] n620_o;
  wire [1:0] n621_o;
  reg [7:0] n622_o;
  wire [1:0] n623_o;
  reg [7:0] n624_o;
  wire n625_o;
  wire [7:0] n626_o;
  wire [7:0] n627_o;
  wire [7:0] n628_o;
  wire [7:0] n629_o;
  wire [7:0] n630_o;
  wire [7:0] n631_o;
  wire [7:0] n632_o;
  wire [7:0] n633_o;
  wire [7:0] n634_o;
  wire [7:0] n635_o;
  wire [7:0] n636_o;
  wire [7:0] n637_o;
  wire [7:0] n638_o;
  wire [7:0] n639_o;
  wire [7:0] n640_o;
  wire [7:0] n641_o;
  wire [7:0] n642_o;
  wire [7:0] n643_o;
  wire [7:0] n644_o;
  wire [7:0] n645_o;
  wire [7:0] n646_o;
  wire [7:0] n647_o;
  wire [7:0] n648_o;
  wire [7:0] n649_o;
  wire [7:0] n650_o;
  wire [7:0] n651_o;
  wire [7:0] n652_o;
  wire [7:0] n653_o;
  wire [7:0] n654_o;
  wire [7:0] n655_o;
  wire [7:0] n656_o;
  wire [7:0] n657_o;
  wire [7:0] n658_o;
  wire [1:0] n659_o;
  reg [7:0] n660_o;
  wire [1:0] n661_o;
  reg [7:0] n662_o;
  wire [1:0] n663_o;
  reg [7:0] n664_o;
  wire [1:0] n665_o;
  reg [7:0] n666_o;
  wire [1:0] n667_o;
  reg [7:0] n668_o;
  wire [1:0] n669_o;
  reg [7:0] n670_o;
  wire [1:0] n671_o;
  reg [7:0] n672_o;
  wire [1:0] n673_o;
  reg [7:0] n674_o;
  wire [1:0] n675_o;
  reg [7:0] n676_o;
  wire [1:0] n677_o;
  reg [7:0] n678_o;
  wire n679_o;
  wire [7:0] n680_o;
  wire n681_o;
  wire n682_o;
  wire n683_o;
  wire n684_o;
  wire n685_o;
  wire n686_o;
  wire n687_o;
  wire n688_o;
  wire n689_o;
  wire n690_o;
  wire n691_o;
  wire n692_o;
  wire n693_o;
  wire n694_o;
  wire n695_o;
  wire n696_o;
  wire n697_o;
  wire n698_o;
  wire n699_o;
  wire n700_o;
  wire n701_o;
  wire n702_o;
  wire n703_o;
  wire n704_o;
  wire n705_o;
  wire n706_o;
  wire n707_o;
  wire n708_o;
  wire n709_o;
  wire n710_o;
  wire n711_o;
  wire n712_o;
  wire n713_o;
  wire n714_o;
  wire n715_o;
  wire n716_o;
  wire n717_o;
  wire n718_o;
  wire n719_o;
  wire n720_o;
  wire n721_o;
  wire n722_o;
  wire n723_o;
  wire n724_o;
  wire n725_o;
  wire n726_o;
  wire n727_o;
  wire n728_o;
  wire n729_o;
  wire n730_o;
  wire n731_o;
  wire n732_o;
  wire n733_o;
  wire n734_o;
  wire n735_o;
  wire n736_o;
  wire n737_o;
  wire n738_o;
  wire n739_o;
  wire n740_o;
  wire n741_o;
  wire n742_o;
  wire n743_o;
  wire n744_o;
  wire n745_o;
  wire n746_o;
  wire n747_o;
  wire n748_o;
  wire n749_o;
  wire n750_o;
  wire [7:0] n751_o;
  wire [7:0] n752_o;
  wire [7:0] n753_o;
  wire [7:0] n754_o;
  wire [7:0] n755_o;
  wire [7:0] n756_o;
  wire [7:0] n757_o;
  wire [7:0] n758_o;
  wire [7:0] n759_o;
  wire [7:0] n760_o;
  wire [7:0] n761_o;
  wire [7:0] n762_o;
  wire [7:0] n763_o;
  wire [7:0] n764_o;
  wire [7:0] n765_o;
  wire [7:0] n766_o;
  wire [7:0] n767_o;
  wire [7:0] n768_o;
  wire [7:0] n769_o;
  wire [7:0] n770_o;
  wire [7:0] n771_o;
  wire [7:0] n772_o;
  wire [7:0] n773_o;
  wire [7:0] n774_o;
  wire [7:0] n775_o;
  wire [7:0] n776_o;
  wire [7:0] n777_o;
  wire [7:0] n778_o;
  wire [7:0] n779_o;
  wire [7:0] n780_o;
  wire [7:0] n781_o;
  wire [7:0] n782_o;
  wire [7:0] n783_o;
  wire [7:0] n784_o;
  wire [7:0] n785_o;
  wire [7:0] n786_o;
  wire [7:0] n787_o;
  wire [7:0] n788_o;
  wire [7:0] n789_o;
  wire [7:0] n790_o;
  wire [7:0] n791_o;
  wire [7:0] n792_o;
  wire [7:0] n793_o;
  wire [7:0] n794_o;
  wire [7:0] n795_o;
  wire [7:0] n796_o;
  wire [7:0] n797_o;
  wire [7:0] n798_o;
  wire [7:0] n799_o;
  wire [7:0] n800_o;
  wire [7:0] n801_o;
  wire [7:0] n802_o;
  wire [7:0] n803_o;
  wire [7:0] n804_o;
  wire [7:0] n805_o;
  wire [7:0] n806_o;
  wire [7:0] n807_o;
  wire [7:0] n808_o;
  wire [7:0] n809_o;
  wire [7:0] n810_o;
  wire [7:0] n811_o;
  wire [7:0] n812_o;
  wire [7:0] n813_o;
  wire [7:0] n814_o;
  wire [255:0] n815_o;
  wire [7:0] n816_o;
  wire [7:0] n817_o;
  wire [7:0] n818_o;
  wire [7:0] n819_o;
  wire [7:0] n820_o;
  wire [7:0] n821_o;
  wire [7:0] n822_o;
  wire [7:0] n823_o;
  wire [7:0] n824_o;
  wire [7:0] n825_o;
  wire [7:0] n826_o;
  wire [7:0] n827_o;
  wire [7:0] n828_o;
  wire [7:0] n829_o;
  wire [7:0] n830_o;
  wire [7:0] n831_o;
  wire [7:0] n832_o;
  wire [7:0] n833_o;
  wire [7:0] n834_o;
  wire [7:0] n835_o;
  wire [7:0] n836_o;
  wire [7:0] n837_o;
  wire [7:0] n838_o;
  wire [7:0] n839_o;
  wire [7:0] n840_o;
  wire [7:0] n841_o;
  wire [7:0] n842_o;
  wire [7:0] n843_o;
  wire [7:0] n844_o;
  wire [7:0] n845_o;
  wire [7:0] n846_o;
  wire [7:0] n847_o;
  wire [1:0] n848_o;
  reg [7:0] n849_o;
  wire [1:0] n850_o;
  reg [7:0] n851_o;
  wire [1:0] n852_o;
  reg [7:0] n853_o;
  wire [1:0] n854_o;
  reg [7:0] n855_o;
  wire [1:0] n856_o;
  reg [7:0] n857_o;
  wire [1:0] n858_o;
  reg [7:0] n859_o;
  wire [1:0] n860_o;
  reg [7:0] n861_o;
  wire [1:0] n862_o;
  reg [7:0] n863_o;
  wire [1:0] n864_o;
  reg [7:0] n865_o;
  wire [1:0] n866_o;
  reg [7:0] n867_o;
  wire n868_o;
  wire [7:0] n869_o;
  wire [7:0] n870_o;
  wire [7:0] n871_o;
  wire [7:0] n872_o;
  wire [7:0] n873_o;
  wire [7:0] n874_o;
  wire [7:0] n875_o;
  wire [7:0] n876_o;
  wire [7:0] n877_o;
  wire [7:0] n878_o;
  wire [7:0] n879_o;
  wire [7:0] n880_o;
  wire [7:0] n881_o;
  wire [7:0] n882_o;
  wire [7:0] n883_o;
  wire [7:0] n884_o;
  wire [7:0] n885_o;
  wire [7:0] n886_o;
  wire [7:0] n887_o;
  wire [7:0] n888_o;
  wire [7:0] n889_o;
  wire [7:0] n890_o;
  wire [7:0] n891_o;
  wire [7:0] n892_o;
  wire [7:0] n893_o;
  wire [7:0] n894_o;
  wire [7:0] n895_o;
  wire [7:0] n896_o;
  wire [7:0] n897_o;
  wire [7:0] n898_o;
  wire [7:0] n899_o;
  wire [7:0] n900_o;
  wire [7:0] n901_o;
  wire [1:0] n902_o;
  reg [7:0] n903_o;
  wire [1:0] n904_o;
  reg [7:0] n905_o;
  wire [1:0] n906_o;
  reg [7:0] n907_o;
  wire [1:0] n908_o;
  reg [7:0] n909_o;
  wire [1:0] n910_o;
  reg [7:0] n911_o;
  wire [1:0] n912_o;
  reg [7:0] n913_o;
  wire [1:0] n914_o;
  reg [7:0] n915_o;
  wire [1:0] n916_o;
  reg [7:0] n917_o;
  wire [1:0] n918_o;
  reg [7:0] n919_o;
  wire [1:0] n920_o;
  reg [7:0] n921_o;
  wire n922_o;
  wire [7:0] n923_o;
  wire n924_o;
  wire n925_o;
  wire n926_o;
  wire n927_o;
  wire n928_o;
  wire n929_o;
  wire n930_o;
  wire n931_o;
  wire n932_o;
  wire n933_o;
  wire n934_o;
  wire n935_o;
  wire n936_o;
  wire n937_o;
  wire n938_o;
  wire n939_o;
  wire n940_o;
  wire n941_o;
  wire n942_o;
  wire n943_o;
  wire n944_o;
  wire n945_o;
  wire n946_o;
  wire n947_o;
  wire n948_o;
  wire n949_o;
  wire n950_o;
  wire n951_o;
  wire n952_o;
  wire n953_o;
  wire n954_o;
  wire n955_o;
  wire n956_o;
  wire n957_o;
  wire n958_o;
  wire n959_o;
  wire n960_o;
  wire n961_o;
  wire n962_o;
  wire n963_o;
  wire n964_o;
  wire n965_o;
  wire n966_o;
  wire n967_o;
  wire n968_o;
  wire n969_o;
  wire n970_o;
  wire n971_o;
  wire n972_o;
  wire n973_o;
  wire n974_o;
  wire n975_o;
  wire n976_o;
  wire n977_o;
  wire n978_o;
  wire n979_o;
  wire n980_o;
  wire n981_o;
  wire n982_o;
  wire n983_o;
  wire n984_o;
  wire n985_o;
  wire n986_o;
  wire n987_o;
  wire n988_o;
  wire n989_o;
  wire n990_o;
  wire n991_o;
  wire n992_o;
  wire n993_o;
  wire [7:0] n994_o;
  wire [7:0] n995_o;
  wire [7:0] n996_o;
  wire [7:0] n997_o;
  wire [7:0] n998_o;
  wire [7:0] n999_o;
  wire [7:0] n1000_o;
  wire [7:0] n1001_o;
  wire [7:0] n1002_o;
  wire [7:0] n1003_o;
  wire [7:0] n1004_o;
  wire [7:0] n1005_o;
  wire [7:0] n1006_o;
  wire [7:0] n1007_o;
  wire [7:0] n1008_o;
  wire [7:0] n1009_o;
  wire [7:0] n1010_o;
  wire [7:0] n1011_o;
  wire [7:0] n1012_o;
  wire [7:0] n1013_o;
  wire [7:0] n1014_o;
  wire [7:0] n1015_o;
  wire [7:0] n1016_o;
  wire [7:0] n1017_o;
  wire [7:0] n1018_o;
  wire [7:0] n1019_o;
  wire [7:0] n1020_o;
  wire [7:0] n1021_o;
  wire [7:0] n1022_o;
  wire [7:0] n1023_o;
  wire [7:0] n1024_o;
  wire [7:0] n1025_o;
  wire [7:0] n1026_o;
  wire [7:0] n1027_o;
  wire [7:0] n1028_o;
  wire [7:0] n1029_o;
  wire [7:0] n1030_o;
  wire [7:0] n1031_o;
  wire [7:0] n1032_o;
  wire [7:0] n1033_o;
  wire [7:0] n1034_o;
  wire [7:0] n1035_o;
  wire [7:0] n1036_o;
  wire [7:0] n1037_o;
  wire [7:0] n1038_o;
  wire [7:0] n1039_o;
  wire [7:0] n1040_o;
  wire [7:0] n1041_o;
  wire [7:0] n1042_o;
  wire [7:0] n1043_o;
  wire [7:0] n1044_o;
  wire [7:0] n1045_o;
  wire [7:0] n1046_o;
  wire [7:0] n1047_o;
  wire [7:0] n1048_o;
  wire [7:0] n1049_o;
  wire [7:0] n1050_o;
  wire [7:0] n1051_o;
  wire [7:0] n1052_o;
  wire [7:0] n1053_o;
  wire [7:0] n1054_o;
  wire [7:0] n1055_o;
  wire [7:0] n1056_o;
  wire [7:0] n1057_o;
  wire [255:0] n1058_o;
  wire [7:0] n1059_o;
  wire [7:0] n1060_o;
  wire [7:0] n1061_o;
  wire [7:0] n1062_o;
  wire [7:0] n1063_o;
  wire [7:0] n1064_o;
  wire [7:0] n1065_o;
  wire [7:0] n1066_o;
  wire [7:0] n1067_o;
  wire [7:0] n1068_o;
  wire [7:0] n1069_o;
  wire [7:0] n1070_o;
  wire [7:0] n1071_o;
  wire [7:0] n1072_o;
  wire [7:0] n1073_o;
  wire [7:0] n1074_o;
  wire [7:0] n1075_o;
  wire [7:0] n1076_o;
  wire [7:0] n1077_o;
  wire [7:0] n1078_o;
  wire [7:0] n1079_o;
  wire [7:0] n1080_o;
  wire [7:0] n1081_o;
  wire [7:0] n1082_o;
  wire [7:0] n1083_o;
  wire [7:0] n1084_o;
  wire [7:0] n1085_o;
  wire [7:0] n1086_o;
  wire [7:0] n1087_o;
  wire [7:0] n1088_o;
  wire [7:0] n1089_o;
  wire [7:0] n1090_o;
  wire [1:0] n1091_o;
  reg [7:0] n1092_o;
  wire [1:0] n1093_o;
  reg [7:0] n1094_o;
  wire [1:0] n1095_o;
  reg [7:0] n1096_o;
  wire [1:0] n1097_o;
  reg [7:0] n1098_o;
  wire [1:0] n1099_o;
  reg [7:0] n1100_o;
  wire [1:0] n1101_o;
  reg [7:0] n1102_o;
  wire [1:0] n1103_o;
  reg [7:0] n1104_o;
  wire [1:0] n1105_o;
  reg [7:0] n1106_o;
  wire [1:0] n1107_o;
  reg [7:0] n1108_o;
  wire [1:0] n1109_o;
  reg [7:0] n1110_o;
  wire n1111_o;
  wire [7:0] n1112_o;
  assign uo_out = n329_o; //(module output)
  assign uio_out = n14_o; //(module output)
  assign uio_oe = n15_o; //(module output)
  /* project.vhdl:21:12  */
  always @*
    rom_mrse = n305_q; // (isignal)
  initial
    rom_mrse = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* project.vhdl:64:12  */
  always @*
    ascell_mrse = n28_o; // (isignal)
  initial
    ascell_mrse = 2'b00;
  /* project.vhdl:65:12  */
  always @*
    cell_mrse = n309_q; // (isignal)
  initial
    cell_mrse = 2'b00;
  /* project.vhdl:66:12  */
  always @*
    ui_in_old = n312_q; // (isignal)
  initial
    ui_in_old = 6'b000000;
  /* project.vhdl:67:12  */
  always @*
    ui_in_sync = n18_o; // (isignal)
  initial
    ui_in_sync = 6'b000000;
  /* project.vhdl:68:12  */
  always @*
    sr_mrse = n315_q; // (isignal)
  initial
    sr_mrse = 8'b00000000;
  /* project.vhdl:69:12  */
  always @*
    i_sr_mrse = n316_q; // (isignal)
  initial
    i_sr_mrse = 3'b000;
  /* project.vhdl:70:12  */
  always @*
    flush_sr_mrse = n320_q; // (isignal)
  initial
    flush_sr_mrse = 1'b0;
  /* project.vhdl:71:12  */
  always @*
    i_rom_mrse = n321_q; // (isignal)
  initial
    i_rom_mrse = 5'b00000;
  /* project.vhdl:73:12  */
  always @*
    time_mrse = n324_q; // (isignal)
  initial
    time_mrse = 14'b00000000000000;
  /* project.vhdl:74:12  */
  always @*
    state_mrse = n327_q; // (isignal)
  initial
    state_mrse = 3'b000;
  /* project.vhdl:80:28  */
  assign n16_o = ui_in[5:0]; // extract
  /* project.vhdl:80:45  */
  assign n17_o = ~ui_in_old;
  /* project.vhdl:80:41  */
  assign n18_o = n16_o & n17_o;
  /* project.vhdl:84:28  */
  assign n21_o = ui_in_sync[0]; // extract
  /* project.vhdl:84:53  */
  assign n22_o = ui_in_sync[1]; // extract
  /* project.vhdl:84:39  */
  assign n23_o = n21_o | n22_o;
  /* project.vhdl:84:70  */
  assign n24_o = ~flush_sr_mrse;
  /* project.vhdl:84:65  */
  assign n25_o = n24_o & n23_o;
  /* project.vhdl:85:42  */
  assign n26_o = ui_in_sync[1:0]; // extract
  /* project.vhdl:84:13  */
  assign n28_o = n25_o ? n26_o : 2'b00;
  /* project.vhdl:137:35  */
  assign n33_o = ui_in[5:0]; // extract
  /* project.vhdl:139:31  */
  assign n35_o = state_mrse == 3'b000;
  /* project.vhdl:140:35  */
  assign n36_o = ui_in_sync[2]; // extract
  /* project.vhdl:140:21  */
  assign n38_o = n36_o ? 1'b1 : flush_sr_mrse;
  /* project.vhdl:144:35  */
  assign n40_o = i_sr_mrse == 3'b100;
  /* project.vhdl:149:50  */
  assign n43_o = {27'b0, i_rom_mrse};  //  uext
  /* project.vhdl:149:50  */
  assign n45_o = n43_o + 32'b00000000000000000000000000000001;
  /* project.vhdl:149:39  */
  assign n46_o = n45_o[4:0];  // trunc
  /* project.vhdl:154:64  */
  assign n47_o = ui_in_sync[0]; // extract
  /* project.vhdl:154:50  */
  assign n48_o = flush_sr_mrse | n47_o;
  /* project.vhdl:154:89  */
  assign n49_o = ui_in_sync[1]; // extract
  /* project.vhdl:154:75  */
  assign n50_o = n48_o | n49_o;
  /* project.vhdl:155:47  */
  assign n51_o = sr_mrse[5:0]; // extract
  /* project.vhdl:155:60  */
  assign n52_o = {n51_o, ascell_mrse};
  /* project.vhdl:157:52  */
  assign n54_o = i_sr_mrse + 3'b001;
  /* project.vhdl:154:21  */
  assign n55_o = n50_o ? n52_o : sr_mrse;
  /* project.vhdl:154:21  */
  assign n56_o = n50_o ? n54_o : i_sr_mrse;
  /* project.vhdl:139:17  */
  assign n57_o = n65_o ? n464_o : rom_mrse;
  /* project.vhdl:144:21  */
  assign n59_o = n40_o ? 8'b00000000 : n55_o;
  /* project.vhdl:144:21  */
  assign n61_o = n40_o ? 3'b000 : n56_o;
  /* project.vhdl:144:21  */
  assign n63_o = n40_o ? 1'b0 : n38_o;
  /* project.vhdl:139:17  */
  assign n64_o = n69_o ? n46_o : i_rom_mrse;
  /* project.vhdl:139:17  */
  assign n65_o = n40_o & n35_o;
  /* project.vhdl:139:17  */
  assign n66_o = n35_o ? n59_o : sr_mrse;
  /* project.vhdl:139:17  */
  assign n67_o = n35_o ? n61_o : i_sr_mrse;
  /* project.vhdl:139:17  */
  assign n69_o = n40_o & n35_o;
  /* project.vhdl:164:30  */
  assign n70_o = ui_in_sync[3]; // extract
  /* project.vhdl:168:33  */
  assign n71_o = ui_in_sync[4]; // extract
  /* project.vhdl:172:33  */
  assign n72_o = ui_in_sync[5]; // extract
  /* project.vhdl:172:17  */
  assign n74_o = n72_o ? 3'b000 : n67_o;
  /* project.vhdl:172:17  */
  assign n76_o = n72_o ? 5'b00000 : n64_o;
  /* project.vhdl:172:17  */
  assign n78_o = n72_o ? 3'b110 : state_mrse;
  /* project.vhdl:168:17  */
  assign n80_o = n71_o ? 3'b000 : n74_o;
  /* project.vhdl:168:17  */
  assign n82_o = n71_o ? 5'b00000 : n76_o;
  /* project.vhdl:168:17  */
  assign n84_o = n71_o ? 3'b101 : n78_o;
  /* project.vhdl:164:17  */
  assign n86_o = n70_o ? 3'b000 : n80_o;
  /* project.vhdl:164:17  */
  assign n88_o = n70_o ? 5'b00000 : n82_o;
  /* project.vhdl:164:17  */
  assign n90_o = n70_o ? 3'b001 : n84_o;
  /* project.vhdl:178:31  */
  assign n92_o = state_mrse == 3'b001;
  /* project.vhdl:179:35  */
  assign n93_o = {27'b0, i_rom_mrse};  //  uext
  /* project.vhdl:179:35  */
  assign n95_o = n93_o == 32'b00000000000000000000000000011111;
  /* project.vhdl:179:21  */
  assign n97_o = n95_o ? 3'b000 : n86_o;
  /* project.vhdl:179:21  */
  assign n99_o = n95_o ? 5'b00000 : n88_o;
  /* project.vhdl:179:21  */
  assign n102_o = n95_o ? 3'b000 : 3'b011;
  /* project.vhdl:187:34  */
  assign n104_o = i_sr_mrse == 3'b011;
  /* project.vhdl:189:50  */
  assign n105_o = {27'b0, i_rom_mrse};  //  uext
  /* project.vhdl:189:50  */
  assign n107_o = n105_o + 32'b00000000000000000000000000000001;
  /* project.vhdl:189:39  */
  assign n108_o = n107_o[4:0];  // trunc
  /* project.vhdl:187:21  */
  assign n110_o = n104_o ? 3'b000 : n97_o;
  /* project.vhdl:187:21  */
  assign n111_o = n104_o ? n108_o : n99_o;
  /* project.vhdl:196:49  */
  assign n114_o = sr_mrse[7:6]; // extract
  /* project.vhdl:195:25  */
  assign n116_o = i_sr_mrse == 3'b000;
  /* project.vhdl:198:49  */
  assign n117_o = sr_mrse[5:4]; // extract
  /* project.vhdl:197:25  */
  assign n119_o = i_sr_mrse == 3'b001;
  /* project.vhdl:200:49  */
  assign n120_o = sr_mrse[3:2]; // extract
  /* project.vhdl:199:25  */
  assign n122_o = i_sr_mrse == 3'b010;
  /* project.vhdl:202:49  */
  assign n123_o = sr_mrse[1:0]; // extract
  /* project.vhdl:201:25  */
  assign n125_o = i_sr_mrse == 3'b011;
  assign n126_o = {n125_o, n122_o, n119_o, n116_o};
  /* project.vhdl:194:21  */
  always @*
    case (n126_o)
      4'b1000: n127_o = n123_o;
      4'b0100: n127_o = n120_o;
      4'b0010: n127_o = n117_o;
      4'b0001: n127_o = n114_o;
      default: n127_o = cell_mrse;
    endcase
  /* project.vhdl:207:34  */
  assign n129_o = state_mrse == 3'b010;
  /* project.vhdl:208:34  */
  assign n130_o = {18'b0, time_mrse};  //  uext
  /* project.vhdl:208:34  */
  assign n132_o = $signed(n130_o) > $signed(32'b00000000000000000000001111101000);
  /* project.vhdl:209:48  */
  assign n133_o = {18'b0, time_mrse};  //  uext
  /* project.vhdl:209:48  */
  assign n135_o = n133_o - 32'b00000000000000000000000000000001;
  /* project.vhdl:209:38  */
  assign n136_o = n135_o[13:0];  // trunc
  /* project.vhdl:211:37  */
  assign n138_o = {18'b0, time_mrse};  //  uext
  /* project.vhdl:211:37  */
  assign n140_o = $signed(n138_o) > $signed(32'b00000000000000000000000000000001);
  /* project.vhdl:213:48  */
  assign n142_o = {18'b0, time_mrse};  //  uext
  /* project.vhdl:213:48  */
  assign n144_o = n142_o - 32'b00000000000000000000000000000001;
  /* project.vhdl:213:38  */
  assign n145_o = n144_o[13:0];  // trunc
  /* project.vhdl:215:48  */
  assign n147_o = i_sr_mrse + 3'b001;
  assign n148_o = n329_o[0]; // extract
  /* project.vhdl:211:21  */
  assign n149_o = n140_o ? 1'b0 : n148_o;
  /* project.vhdl:211:21  */
  assign n150_o = n140_o ? n86_o : n147_o;
  /* project.vhdl:211:21  */
  assign n151_o = n140_o ? n145_o : time_mrse;
  /* project.vhdl:211:21  */
  assign n153_o = n140_o ? n90_o : 3'b001;
  /* project.vhdl:208:21  */
  assign n154_o = n132_o ? 1'b1 : n149_o;
  /* project.vhdl:208:21  */
  assign n155_o = n132_o ? n86_o : n150_o;
  /* project.vhdl:208:21  */
  assign n156_o = n132_o ? n136_o : n151_o;
  /* project.vhdl:208:21  */
  assign n157_o = n132_o ? n90_o : n153_o;
  /* project.vhdl:218:34  */
  assign n159_o = state_mrse == 3'b011;
  /* project.vhdl:223:40  */
  assign n163_o = sr_mrse == 8'b00000000;
  /* project.vhdl:224:56  */
  assign n165_o = i_sr_mrse + 3'b001;
  /* project.vhdl:223:29  */
  assign n166_o = n163_o ? n165_o : n86_o;
  /* project.vhdl:220:25  */
  assign n168_o = cell_mrse == 2'b00;
  /* project.vhdl:230:40  */
  assign n172_o = sr_mrse == 8'b11111111;
  /* project.vhdl:231:56  */
  assign n174_o = i_sr_mrse + 3'b001;
  /* project.vhdl:230:29  */
  assign n175_o = n172_o ? n174_o : n86_o;
  /* project.vhdl:227:25  */
  assign n177_o = cell_mrse == 2'b11;
  /* project.vhdl:234:25  */
  assign n179_o = cell_mrse == 2'b01;
  /* project.vhdl:237:25  */
  assign n181_o = cell_mrse == 2'b10;
  assign n182_o = {n181_o, n179_o, n177_o, n168_o};
  /* project.vhdl:219:21  */
  always @*
    case (n182_o)
      4'b1000: n183_o = n66_o;
      4'b0100: n183_o = n66_o;
      4'b0010: n183_o = n626_o;
      4'b0001: n183_o = n572_o;
      default: n183_o = n66_o;
    endcase
  /* project.vhdl:219:21  */
  always @*
    case (n182_o)
      4'b1000: n184_o = n86_o;
      4'b0100: n184_o = n86_o;
      4'b0010: n184_o = n175_o;
      4'b0001: n184_o = n166_o;
      default: n184_o = n86_o;
    endcase
  /* project.vhdl:219:21  */
  always @*
    case (n182_o)
      4'b1000: n187_o = 14'b01011101110000;
      4'b0100: n187_o = 14'b00101110111000;
      4'b0010: n187_o = time_mrse;
      4'b0001: n187_o = time_mrse;
      default: n187_o = time_mrse;
    endcase
  /* project.vhdl:219:21  */
  always @*
    case (n182_o)
      4'b1000: n192_o = 3'b010;
      4'b0100: n192_o = 3'b010;
      4'b0010: n192_o = 3'b001;
      4'b0001: n192_o = 3'b001;
      default: n192_o = n90_o;
    endcase
  /* project.vhdl:244:34  */
  assign n194_o = state_mrse == 3'b101;
  /* project.vhdl:245:35  */
  assign n195_o = {27'b0, i_rom_mrse};  //  uext
  /* project.vhdl:245:35  */
  assign n197_o = $signed(n195_o) < $signed(32'b00000000000000000000000000011111);
  /* project.vhdl:246:36  */
  assign n200_o = sr_mrse == n680_o;
  /* project.vhdl:247:53  */
  assign n202_o = ~sr_mrse;
  /* project.vhdl:248:54  */
  assign n204_o = {27'b0, i_rom_mrse};  //  uext
  /* project.vhdl:248:54  */
  assign n206_o = n204_o + 32'b00000000000000000000000000000001;
  /* project.vhdl:248:43  */
  assign n207_o = n206_o[4:0];  // trunc
  /* project.vhdl:245:21  */
  assign n210_o = n213_o ? n815_o : n57_o;
  /* project.vhdl:246:25  */
  assign n211_o = n200_o ? n66_o : n869_o;
  /* project.vhdl:246:25  */
  assign n212_o = n200_o ? n207_o : n88_o;
  /* project.vhdl:245:21  */
  assign n213_o = n200_o & n197_o;
  /* project.vhdl:245:21  */
  assign n214_o = n197_o ? n211_o : n66_o;
  /* project.vhdl:245:21  */
  assign n216_o = n197_o ? n212_o : 5'b00000;
  /* project.vhdl:245:21  */
  assign n218_o = n197_o ? n90_o : 3'b000;
  /* project.vhdl:257:34  */
  assign n220_o = state_mrse == 3'b110;
  /* project.vhdl:258:35  */
  assign n221_o = {27'b0, i_rom_mrse};  //  uext
  /* project.vhdl:258:35  */
  assign n223_o = $signed(n221_o) < $signed(32'b00000000000000000000000000011111);
  /* project.vhdl:259:36  */
  assign n226_o = sr_mrse == n923_o;
  /* project.vhdl:260:53  */
  assign n228_o = ~sr_mrse;
  /* project.vhdl:261:54  */
  assign n230_o = {27'b0, i_rom_mrse};  //  uext
  /* project.vhdl:261:54  */
  assign n232_o = n230_o + 32'b00000000000000000000000000000001;
  /* project.vhdl:261:43  */
  assign n233_o = n232_o[4:0];  // trunc
  /* project.vhdl:257:17  */
  assign n236_o = n245_o ? n1058_o : n57_o;
  /* project.vhdl:259:25  */
  assign n237_o = n226_o ? n66_o : n1112_o;
  /* project.vhdl:259:25  */
  assign n238_o = n226_o ? n233_o : n88_o;
  /* project.vhdl:258:21  */
  assign n239_o = n226_o & n223_o;
  /* project.vhdl:257:17  */
  assign n240_o = n246_o ? n237_o : n66_o;
  /* project.vhdl:258:21  */
  assign n242_o = n223_o ? n238_o : 5'b00000;
  /* project.vhdl:258:21  */
  assign n244_o = n223_o ? n90_o : 3'b000;
  /* project.vhdl:257:17  */
  assign n245_o = n239_o & n220_o;
  /* project.vhdl:257:17  */
  assign n246_o = n223_o & n220_o;
  /* project.vhdl:257:17  */
  assign n247_o = n220_o ? n242_o : n88_o;
  /* project.vhdl:257:17  */
  assign n248_o = n220_o ? n244_o : n90_o;
  /* project.vhdl:244:17  */
  assign n249_o = n194_o ? n210_o : n236_o;
  /* project.vhdl:244:17  */
  assign n250_o = n194_o ? n214_o : n240_o;
  /* project.vhdl:244:17  */
  assign n251_o = n194_o ? n216_o : n247_o;
  /* project.vhdl:244:17  */
  assign n252_o = n194_o ? n218_o : n248_o;
  /* project.vhdl:218:17  */
  assign n253_o = n159_o ? n57_o : n249_o;
  /* project.vhdl:218:17  */
  assign n254_o = n159_o ? n183_o : n250_o;
  /* project.vhdl:218:17  */
  assign n255_o = n159_o ? n184_o : n86_o;
  /* project.vhdl:218:17  */
  assign n256_o = n159_o ? n88_o : n251_o;
  /* project.vhdl:218:17  */
  assign n257_o = n159_o ? n187_o : time_mrse;
  /* project.vhdl:218:17  */
  assign n258_o = n159_o ? n192_o : n252_o;
  assign n259_o = n329_o[0]; // extract
  /* project.vhdl:207:17  */
  assign n260_o = n129_o ? n154_o : n259_o;
  /* project.vhdl:207:17  */
  assign n261_o = n129_o ? n57_o : n253_o;
  /* project.vhdl:207:17  */
  assign n262_o = n129_o ? n66_o : n254_o;
  /* project.vhdl:207:17  */
  assign n263_o = n129_o ? n155_o : n255_o;
  /* project.vhdl:207:17  */
  assign n264_o = n129_o ? n88_o : n256_o;
  /* project.vhdl:207:17  */
  assign n265_o = n129_o ? n156_o : n257_o;
  /* project.vhdl:207:17  */
  assign n266_o = n129_o ? n157_o : n258_o;
  assign n267_o = n329_o[0]; // extract
  /* project.vhdl:178:17  */
  assign n268_o = n92_o ? n267_o : n260_o;
  /* project.vhdl:178:17  */
  assign n269_o = n92_o ? n57_o : n261_o;
  /* project.vhdl:178:17  */
  assign n271_o = n92_o ? n518_o : n262_o;
  /* project.vhdl:178:17  */
  assign n272_o = n92_o ? n110_o : n263_o;
  /* project.vhdl:178:17  */
  assign n273_o = n92_o ? n111_o : n264_o;
  /* project.vhdl:178:17  */
  assign n274_o = n92_o ? time_mrse : n265_o;
  /* project.vhdl:178:17  */
  assign n275_o = n92_o ? n102_o : n266_o;
  assign n290_o = n329_o[7:1]; // extract
  /* project.vhdl:95:13  */
  assign n291_o = rst_n ? 7'b0000000 : n290_o;
  /* project.vhdl:135:13  */
  always @(posedge clk or posedge rst_n)
    if (rst_n)
      n305_q <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n305_q <= n269_o;
  /* project.vhdl:92:9  */
  assign n306_o = ~rst_n;
  /* project.vhdl:92:9  */
  assign n307_o = n92_o & n306_o;
  /* project.vhdl:135:13  */
  assign n308_o = n307_o ? n127_o : cell_mrse;
  /* project.vhdl:135:13  */
  always @(posedge clk)
    n309_q <= n308_o;
  initial
    n309_q = 2'b00;
  /* project.vhdl:92:9  */
  assign n310_o = ~rst_n;
  /* project.vhdl:135:13  */
  assign n311_o = n310_o ? n33_o : ui_in_old;
  /* project.vhdl:135:13  */
  always @(posedge clk)
    n312_q <= n311_o;
  initial
    n312_q = 6'b000000;
  /* project.vhdl:92:9  */
  assign n313_o = ~rst_n;
  /* project.vhdl:135:13  */
  assign n314_o = n313_o ? n271_o : sr_mrse;
  /* project.vhdl:135:13  */
  always @(posedge clk)
    n315_q <= n314_o;
  initial
    n315_q = 8'b00000000;
  /* project.vhdl:135:13  */
  always @(posedge clk or posedge rst_n)
    if (rst_n)
      n316_q <= 3'b000;
    else
      n316_q <= n272_o;
  /* project.vhdl:92:9  */
  assign n317_o = ~rst_n;
  /* project.vhdl:92:9  */
  assign n318_o = n35_o & n317_o;
  /* project.vhdl:135:13  */
  assign n319_o = n318_o ? n63_o : flush_sr_mrse;
  /* project.vhdl:135:13  */
  always @(posedge clk)
    n320_q <= n319_o;
  initial
    n320_q = 1'b0;
  /* project.vhdl:135:13  */
  always @(posedge clk or posedge rst_n)
    if (rst_n)
      n321_q <= 5'b00000;
    else
      n321_q <= n273_o;
  /* project.vhdl:92:9  */
  assign n322_o = ~rst_n;
  /* project.vhdl:135:13  */
  assign n323_o = n322_o ? n274_o : time_mrse;
  /* project.vhdl:135:13  */
  always @(posedge clk)
    n324_q <= n323_o;
  initial
    n324_q = 14'b00000000000000;
  /* project.vhdl:92:9  */
  assign n325_o = ~rst_n;
  /* project.vhdl:135:13  */
  assign n326_o = n325_o ? n275_o : state_mrse;
  /* project.vhdl:135:13  */
  always @(posedge clk)
    n327_q <= n326_o;
  initial
    n327_q = 3'b000;
  /* project.vhdl:135:13  */
  always @(posedge clk or posedge rst_n)
    if (rst_n)
      n328_q <= 1'b0;
    else
      n328_q <= n268_o;
  /* project.vhdl:95:13  */
  assign n329_o = {n291_o, n328_q};
  /* project.vhdl:148:25  */
  assign n330_o = i_rom_mrse[4]; // extract
  /* project.vhdl:148:25  */
  assign n331_o = ~n330_o;
  /* project.vhdl:148:25  */
  assign n332_o = i_rom_mrse[3]; // extract
  /* project.vhdl:148:25  */
  assign n333_o = ~n332_o;
  /* project.vhdl:148:25  */
  assign n334_o = n331_o & n333_o;
  /* project.vhdl:148:25  */
  assign n335_o = n331_o & n332_o;
  /* project.vhdl:148:25  */
  assign n336_o = n330_o & n333_o;
  /* project.vhdl:148:25  */
  assign n337_o = n330_o & n332_o;
  /* project.vhdl:148:25  */
  assign n338_o = i_rom_mrse[2]; // extract
  /* project.vhdl:148:25  */
  assign n339_o = ~n338_o;
  /* project.vhdl:148:25  */
  assign n340_o = n334_o & n339_o;
  /* project.vhdl:148:25  */
  assign n341_o = n334_o & n338_o;
  /* project.vhdl:148:25  */
  assign n342_o = n335_o & n339_o;
  /* project.vhdl:148:25  */
  assign n343_o = n335_o & n338_o;
  /* project.vhdl:148:25  */
  assign n344_o = n336_o & n339_o;
  /* project.vhdl:148:25  */
  assign n345_o = n336_o & n338_o;
  /* project.vhdl:148:25  */
  assign n346_o = n337_o & n339_o;
  /* project.vhdl:148:25  */
  assign n347_o = n337_o & n338_o;
  /* project.vhdl:148:25  */
  assign n348_o = i_rom_mrse[1]; // extract
  /* project.vhdl:148:25  */
  assign n349_o = ~n348_o;
  /* project.vhdl:148:25  */
  assign n350_o = n340_o & n349_o;
  /* project.vhdl:148:25  */
  assign n351_o = n340_o & n348_o;
  /* project.vhdl:148:25  */
  assign n352_o = n341_o & n349_o;
  /* project.vhdl:148:25  */
  assign n353_o = n341_o & n348_o;
  /* project.vhdl:148:25  */
  assign n354_o = n342_o & n349_o;
  /* project.vhdl:148:25  */
  assign n355_o = n342_o & n348_o;
  /* project.vhdl:148:25  */
  assign n356_o = n343_o & n349_o;
  /* project.vhdl:148:25  */
  assign n357_o = n343_o & n348_o;
  /* project.vhdl:148:25  */
  assign n358_o = n344_o & n349_o;
  /* project.vhdl:148:25  */
  assign n359_o = n344_o & n348_o;
  /* project.vhdl:148:25  */
  assign n360_o = n345_o & n349_o;
  /* project.vhdl:148:25  */
  assign n361_o = n345_o & n348_o;
  /* project.vhdl:148:25  */
  assign n362_o = n346_o & n349_o;
  /* project.vhdl:148:25  */
  assign n363_o = n346_o & n348_o;
  /* project.vhdl:148:25  */
  assign n364_o = n347_o & n349_o;
  /* project.vhdl:148:25  */
  assign n365_o = n347_o & n348_o;
  /* project.vhdl:148:25  */
  assign n366_o = i_rom_mrse[0]; // extract
  /* project.vhdl:148:25  */
  assign n367_o = ~n366_o;
  /* project.vhdl:148:25  */
  assign n368_o = n350_o & n367_o;
  /* project.vhdl:148:25  */
  assign n369_o = n350_o & n366_o;
  /* project.vhdl:148:25  */
  assign n370_o = n351_o & n367_o;
  /* project.vhdl:148:25  */
  assign n371_o = n351_o & n366_o;
  /* project.vhdl:148:25  */
  assign n372_o = n352_o & n367_o;
  /* project.vhdl:148:25  */
  assign n373_o = n352_o & n366_o;
  /* project.vhdl:148:25  */
  assign n374_o = n353_o & n367_o;
  /* project.vhdl:148:25  */
  assign n375_o = n353_o & n366_o;
  /* project.vhdl:148:25  */
  assign n376_o = n354_o & n367_o;
  /* project.vhdl:148:25  */
  assign n377_o = n354_o & n366_o;
  /* project.vhdl:148:25  */
  assign n378_o = n355_o & n367_o;
  /* project.vhdl:148:25  */
  assign n379_o = n355_o & n366_o;
  /* project.vhdl:148:25  */
  assign n380_o = n356_o & n367_o;
  /* project.vhdl:148:25  */
  assign n381_o = n356_o & n366_o;
  /* project.vhdl:148:25  */
  assign n382_o = n357_o & n367_o;
  /* project.vhdl:148:25  */
  assign n383_o = n357_o & n366_o;
  /* project.vhdl:148:25  */
  assign n384_o = n358_o & n367_o;
  /* project.vhdl:148:25  */
  assign n385_o = n358_o & n366_o;
  /* project.vhdl:148:25  */
  assign n386_o = n359_o & n367_o;
  /* project.vhdl:148:25  */
  assign n387_o = n359_o & n366_o;
  /* project.vhdl:148:25  */
  assign n388_o = n360_o & n367_o;
  /* project.vhdl:148:25  */
  assign n389_o = n360_o & n366_o;
  /* project.vhdl:148:25  */
  assign n390_o = n361_o & n367_o;
  /* project.vhdl:148:25  */
  assign n391_o = n361_o & n366_o;
  /* project.vhdl:148:25  */
  assign n392_o = n362_o & n367_o;
  /* project.vhdl:148:25  */
  assign n393_o = n362_o & n366_o;
  /* project.vhdl:148:25  */
  assign n394_o = n363_o & n367_o;
  /* project.vhdl:148:25  */
  assign n395_o = n363_o & n366_o;
  /* project.vhdl:148:25  */
  assign n396_o = n364_o & n367_o;
  /* project.vhdl:148:25  */
  assign n397_o = n364_o & n366_o;
  /* project.vhdl:148:25  */
  assign n398_o = n365_o & n367_o;
  /* project.vhdl:148:25  */
  assign n399_o = n365_o & n366_o;
  assign n400_o = rom_mrse[7:0]; // extract
  /* project.vhdl:148:25  */
  assign n401_o = n368_o ? sr_mrse : n400_o;
  assign n402_o = rom_mrse[15:8]; // extract
  /* project.vhdl:148:25  */
  assign n403_o = n369_o ? sr_mrse : n402_o;
  assign n404_o = rom_mrse[23:16]; // extract
  /* project.vhdl:148:25  */
  assign n405_o = n370_o ? sr_mrse : n404_o;
  assign n406_o = rom_mrse[31:24]; // extract
  /* project.vhdl:148:25  */
  assign n407_o = n371_o ? sr_mrse : n406_o;
  assign n408_o = rom_mrse[39:32]; // extract
  /* project.vhdl:148:25  */
  assign n409_o = n372_o ? sr_mrse : n408_o;
  assign n410_o = rom_mrse[47:40]; // extract
  /* project.vhdl:148:25  */
  assign n411_o = n373_o ? sr_mrse : n410_o;
  assign n412_o = rom_mrse[55:48]; // extract
  /* project.vhdl:148:25  */
  assign n413_o = n374_o ? sr_mrse : n412_o;
  assign n414_o = rom_mrse[63:56]; // extract
  /* project.vhdl:148:25  */
  assign n415_o = n375_o ? sr_mrse : n414_o;
  assign n416_o = rom_mrse[71:64]; // extract
  /* project.vhdl:148:25  */
  assign n417_o = n376_o ? sr_mrse : n416_o;
  assign n418_o = rom_mrse[79:72]; // extract
  /* project.vhdl:148:25  */
  assign n419_o = n377_o ? sr_mrse : n418_o;
  assign n420_o = rom_mrse[87:80]; // extract
  /* project.vhdl:148:25  */
  assign n421_o = n378_o ? sr_mrse : n420_o;
  assign n422_o = rom_mrse[95:88]; // extract
  /* project.vhdl:148:25  */
  assign n423_o = n379_o ? sr_mrse : n422_o;
  assign n424_o = rom_mrse[103:96]; // extract
  /* project.vhdl:148:25  */
  assign n425_o = n380_o ? sr_mrse : n424_o;
  assign n426_o = rom_mrse[111:104]; // extract
  /* project.vhdl:148:25  */
  assign n427_o = n381_o ? sr_mrse : n426_o;
  assign n428_o = rom_mrse[119:112]; // extract
  /* project.vhdl:148:25  */
  assign n429_o = n382_o ? sr_mrse : n428_o;
  assign n430_o = rom_mrse[127:120]; // extract
  /* project.vhdl:148:25  */
  assign n431_o = n383_o ? sr_mrse : n430_o;
  assign n432_o = rom_mrse[135:128]; // extract
  /* project.vhdl:148:25  */
  assign n433_o = n384_o ? sr_mrse : n432_o;
  assign n434_o = rom_mrse[143:136]; // extract
  /* project.vhdl:148:25  */
  assign n435_o = n385_o ? sr_mrse : n434_o;
  assign n436_o = rom_mrse[151:144]; // extract
  /* project.vhdl:148:25  */
  assign n437_o = n386_o ? sr_mrse : n436_o;
  assign n438_o = rom_mrse[159:152]; // extract
  /* project.vhdl:148:25  */
  assign n439_o = n387_o ? sr_mrse : n438_o;
  assign n440_o = rom_mrse[167:160]; // extract
  /* project.vhdl:148:25  */
  assign n441_o = n388_o ? sr_mrse : n440_o;
  assign n442_o = rom_mrse[175:168]; // extract
  /* project.vhdl:148:25  */
  assign n443_o = n389_o ? sr_mrse : n442_o;
  assign n444_o = rom_mrse[183:176]; // extract
  /* project.vhdl:148:25  */
  assign n445_o = n390_o ? sr_mrse : n444_o;
  assign n446_o = rom_mrse[191:184]; // extract
  /* project.vhdl:148:25  */
  assign n447_o = n391_o ? sr_mrse : n446_o;
  assign n448_o = rom_mrse[199:192]; // extract
  /* project.vhdl:148:25  */
  assign n449_o = n392_o ? sr_mrse : n448_o;
  assign n450_o = rom_mrse[207:200]; // extract
  /* project.vhdl:148:25  */
  assign n451_o = n393_o ? sr_mrse : n450_o;
  assign n452_o = rom_mrse[215:208]; // extract
  /* project.vhdl:148:25  */
  assign n453_o = n394_o ? sr_mrse : n452_o;
  assign n454_o = rom_mrse[223:216]; // extract
  /* project.vhdl:148:25  */
  assign n455_o = n395_o ? sr_mrse : n454_o;
  assign n456_o = rom_mrse[231:224]; // extract
  /* project.vhdl:148:25  */
  assign n457_o = n396_o ? sr_mrse : n456_o;
  assign n458_o = rom_mrse[239:232]; // extract
  /* project.vhdl:148:25  */
  assign n459_o = n397_o ? sr_mrse : n458_o;
  assign n460_o = rom_mrse[247:240]; // extract
  /* project.vhdl:148:25  */
  assign n461_o = n398_o ? sr_mrse : n460_o;
  assign n462_o = rom_mrse[255:248]; // extract
  /* project.vhdl:148:25  */
  assign n463_o = n399_o ? sr_mrse : n462_o;
  assign n464_o = {n463_o, n461_o, n459_o, n457_o, n455_o, n453_o, n451_o, n449_o, n447_o, n445_o, n443_o, n441_o, n439_o, n437_o, n435_o, n433_o, n431_o, n429_o, n427_o, n425_o, n423_o, n421_o, n419_o, n417_o, n415_o, n413_o, n411_o, n409_o, n407_o, n405_o, n403_o, n401_o};
  /* project.vhdl:148:34  */
  assign n465_o = rom_mrse[7:0]; // extract
  /* project.vhdl:148:25  */
  assign n466_o = rom_mrse[15:8]; // extract
  assign n467_o = rom_mrse[23:16]; // extract
  assign n468_o = rom_mrse[31:24]; // extract
  assign n469_o = rom_mrse[39:32]; // extract
  assign n470_o = rom_mrse[47:40]; // extract
  assign n471_o = rom_mrse[55:48]; // extract
  assign n472_o = rom_mrse[63:56]; // extract
  assign n473_o = rom_mrse[71:64]; // extract
  assign n474_o = rom_mrse[79:72]; // extract
  assign n475_o = rom_mrse[87:80]; // extract
  assign n476_o = rom_mrse[95:88]; // extract
  assign n477_o = rom_mrse[103:96]; // extract
  assign n478_o = rom_mrse[111:104]; // extract
  assign n479_o = rom_mrse[119:112]; // extract
  assign n480_o = rom_mrse[127:120]; // extract
  assign n481_o = rom_mrse[135:128]; // extract
  assign n482_o = rom_mrse[143:136]; // extract
  assign n483_o = rom_mrse[151:144]; // extract
  assign n484_o = rom_mrse[159:152]; // extract
  assign n485_o = rom_mrse[167:160]; // extract
  assign n486_o = rom_mrse[175:168]; // extract
  assign n487_o = rom_mrse[183:176]; // extract
  assign n488_o = rom_mrse[191:184]; // extract
  assign n489_o = rom_mrse[199:192]; // extract
  assign n490_o = rom_mrse[207:200]; // extract
  assign n491_o = rom_mrse[215:208]; // extract
  assign n492_o = rom_mrse[223:216]; // extract
  assign n493_o = rom_mrse[231:224]; // extract
  assign n494_o = rom_mrse[239:232]; // extract
  assign n495_o = rom_mrse[247:240]; // extract
  assign n496_o = rom_mrse[255:248]; // extract
  /* project.vhdl:192:40  */
  assign n497_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n497_o)
      2'b00: n498_o = n465_o;
      2'b01: n498_o = n466_o;
      2'b10: n498_o = n467_o;
      2'b11: n498_o = n468_o;
    endcase
  /* project.vhdl:192:40  */
  assign n499_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n499_o)
      2'b00: n500_o = n469_o;
      2'b01: n500_o = n470_o;
      2'b10: n500_o = n471_o;
      2'b11: n500_o = n472_o;
    endcase
  /* project.vhdl:192:40  */
  assign n501_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n501_o)
      2'b00: n502_o = n473_o;
      2'b01: n502_o = n474_o;
      2'b10: n502_o = n475_o;
      2'b11: n502_o = n476_o;
    endcase
  /* project.vhdl:192:40  */
  assign n503_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n503_o)
      2'b00: n504_o = n477_o;
      2'b01: n504_o = n478_o;
      2'b10: n504_o = n479_o;
      2'b11: n504_o = n480_o;
    endcase
  /* project.vhdl:192:40  */
  assign n505_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n505_o)
      2'b00: n506_o = n481_o;
      2'b01: n506_o = n482_o;
      2'b10: n506_o = n483_o;
      2'b11: n506_o = n484_o;
    endcase
  /* project.vhdl:192:40  */
  assign n507_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n507_o)
      2'b00: n508_o = n485_o;
      2'b01: n508_o = n486_o;
      2'b10: n508_o = n487_o;
      2'b11: n508_o = n488_o;
    endcase
  /* project.vhdl:192:40  */
  assign n509_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n509_o)
      2'b00: n510_o = n489_o;
      2'b01: n510_o = n490_o;
      2'b10: n510_o = n491_o;
      2'b11: n510_o = n492_o;
    endcase
  /* project.vhdl:192:40  */
  assign n511_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n511_o)
      2'b00: n512_o = n493_o;
      2'b01: n512_o = n494_o;
      2'b10: n512_o = n495_o;
      2'b11: n512_o = n496_o;
    endcase
  /* project.vhdl:192:40  */
  assign n513_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n513_o)
      2'b00: n514_o = n498_o;
      2'b01: n514_o = n500_o;
      2'b10: n514_o = n502_o;
      2'b11: n514_o = n504_o;
    endcase
  /* project.vhdl:192:40  */
  assign n515_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:192:40  */
  always @*
    case (n515_o)
      2'b00: n516_o = n506_o;
      2'b01: n516_o = n508_o;
      2'b10: n516_o = n510_o;
      2'b11: n516_o = n512_o;
    endcase
  /* project.vhdl:192:40  */
  assign n517_o = i_rom_mrse[4]; // extract
  /* project.vhdl:192:40  */
  assign n518_o = n517_o ? n516_o : n514_o;
  /* project.vhdl:192:40  */
  assign n519_o = rom_mrse[7:0]; // extract
  /* project.vhdl:192:41  */
  assign n520_o = rom_mrse[15:8]; // extract
  assign n521_o = rom_mrse[23:16]; // extract
  assign n522_o = rom_mrse[31:24]; // extract
  assign n523_o = rom_mrse[39:32]; // extract
  assign n524_o = rom_mrse[47:40]; // extract
  assign n525_o = rom_mrse[55:48]; // extract
  assign n526_o = rom_mrse[63:56]; // extract
  assign n527_o = rom_mrse[71:64]; // extract
  assign n528_o = rom_mrse[79:72]; // extract
  assign n529_o = rom_mrse[87:80]; // extract
  assign n530_o = rom_mrse[95:88]; // extract
  assign n531_o = rom_mrse[103:96]; // extract
  assign n532_o = rom_mrse[111:104]; // extract
  assign n533_o = rom_mrse[119:112]; // extract
  assign n534_o = rom_mrse[127:120]; // extract
  assign n535_o = rom_mrse[135:128]; // extract
  assign n536_o = rom_mrse[143:136]; // extract
  assign n537_o = rom_mrse[151:144]; // extract
  assign n538_o = rom_mrse[159:152]; // extract
  assign n539_o = rom_mrse[167:160]; // extract
  assign n540_o = rom_mrse[175:168]; // extract
  assign n541_o = rom_mrse[183:176]; // extract
  assign n542_o = rom_mrse[191:184]; // extract
  assign n543_o = rom_mrse[199:192]; // extract
  assign n544_o = rom_mrse[207:200]; // extract
  assign n545_o = rom_mrse[215:208]; // extract
  assign n546_o = rom_mrse[223:216]; // extract
  assign n547_o = rom_mrse[231:224]; // extract
  assign n548_o = rom_mrse[239:232]; // extract
  assign n549_o = rom_mrse[247:240]; // extract
  assign n550_o = rom_mrse[255:248]; // extract
  /* project.vhdl:221:48  */
  assign n551_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n551_o)
      2'b00: n552_o = n519_o;
      2'b01: n552_o = n520_o;
      2'b10: n552_o = n521_o;
      2'b11: n552_o = n522_o;
    endcase
  /* project.vhdl:221:48  */
  assign n553_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n553_o)
      2'b00: n554_o = n523_o;
      2'b01: n554_o = n524_o;
      2'b10: n554_o = n525_o;
      2'b11: n554_o = n526_o;
    endcase
  /* project.vhdl:221:48  */
  assign n555_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n555_o)
      2'b00: n556_o = n527_o;
      2'b01: n556_o = n528_o;
      2'b10: n556_o = n529_o;
      2'b11: n556_o = n530_o;
    endcase
  /* project.vhdl:221:48  */
  assign n557_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n557_o)
      2'b00: n558_o = n531_o;
      2'b01: n558_o = n532_o;
      2'b10: n558_o = n533_o;
      2'b11: n558_o = n534_o;
    endcase
  /* project.vhdl:221:48  */
  assign n559_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n559_o)
      2'b00: n560_o = n535_o;
      2'b01: n560_o = n536_o;
      2'b10: n560_o = n537_o;
      2'b11: n560_o = n538_o;
    endcase
  /* project.vhdl:221:48  */
  assign n561_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n561_o)
      2'b00: n562_o = n539_o;
      2'b01: n562_o = n540_o;
      2'b10: n562_o = n541_o;
      2'b11: n562_o = n542_o;
    endcase
  /* project.vhdl:221:48  */
  assign n563_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n563_o)
      2'b00: n564_o = n543_o;
      2'b01: n564_o = n544_o;
      2'b10: n564_o = n545_o;
      2'b11: n564_o = n546_o;
    endcase
  /* project.vhdl:221:48  */
  assign n565_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n565_o)
      2'b00: n566_o = n547_o;
      2'b01: n566_o = n548_o;
      2'b10: n566_o = n549_o;
      2'b11: n566_o = n550_o;
    endcase
  /* project.vhdl:221:48  */
  assign n567_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n567_o)
      2'b00: n568_o = n552_o;
      2'b01: n568_o = n554_o;
      2'b10: n568_o = n556_o;
      2'b11: n568_o = n558_o;
    endcase
  /* project.vhdl:221:48  */
  assign n569_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:221:48  */
  always @*
    case (n569_o)
      2'b00: n570_o = n560_o;
      2'b01: n570_o = n562_o;
      2'b10: n570_o = n564_o;
      2'b11: n570_o = n566_o;
    endcase
  /* project.vhdl:221:48  */
  assign n571_o = i_rom_mrse[4]; // extract
  /* project.vhdl:221:48  */
  assign n572_o = n571_o ? n570_o : n568_o;
  /* project.vhdl:221:48  */
  assign n573_o = rom_mrse[7:0]; // extract
  /* project.vhdl:221:49  */
  assign n574_o = rom_mrse[15:8]; // extract
  assign n575_o = rom_mrse[23:16]; // extract
  assign n576_o = rom_mrse[31:24]; // extract
  assign n577_o = rom_mrse[39:32]; // extract
  assign n578_o = rom_mrse[47:40]; // extract
  assign n579_o = rom_mrse[55:48]; // extract
  assign n580_o = rom_mrse[63:56]; // extract
  assign n581_o = rom_mrse[71:64]; // extract
  assign n582_o = rom_mrse[79:72]; // extract
  assign n583_o = rom_mrse[87:80]; // extract
  assign n584_o = rom_mrse[95:88]; // extract
  assign n585_o = rom_mrse[103:96]; // extract
  assign n586_o = rom_mrse[111:104]; // extract
  assign n587_o = rom_mrse[119:112]; // extract
  assign n588_o = rom_mrse[127:120]; // extract
  assign n589_o = rom_mrse[135:128]; // extract
  assign n590_o = rom_mrse[143:136]; // extract
  assign n591_o = rom_mrse[151:144]; // extract
  assign n592_o = rom_mrse[159:152]; // extract
  assign n593_o = rom_mrse[167:160]; // extract
  assign n594_o = rom_mrse[175:168]; // extract
  assign n595_o = rom_mrse[183:176]; // extract
  assign n596_o = rom_mrse[191:184]; // extract
  assign n597_o = rom_mrse[199:192]; // extract
  assign n598_o = rom_mrse[207:200]; // extract
  assign n599_o = rom_mrse[215:208]; // extract
  assign n600_o = rom_mrse[223:216]; // extract
  assign n601_o = rom_mrse[231:224]; // extract
  assign n602_o = rom_mrse[239:232]; // extract
  assign n603_o = rom_mrse[247:240]; // extract
  assign n604_o = rom_mrse[255:248]; // extract
  /* project.vhdl:228:48  */
  assign n605_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n605_o)
      2'b00: n606_o = n573_o;
      2'b01: n606_o = n574_o;
      2'b10: n606_o = n575_o;
      2'b11: n606_o = n576_o;
    endcase
  /* project.vhdl:228:48  */
  assign n607_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n607_o)
      2'b00: n608_o = n577_o;
      2'b01: n608_o = n578_o;
      2'b10: n608_o = n579_o;
      2'b11: n608_o = n580_o;
    endcase
  /* project.vhdl:228:48  */
  assign n609_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n609_o)
      2'b00: n610_o = n581_o;
      2'b01: n610_o = n582_o;
      2'b10: n610_o = n583_o;
      2'b11: n610_o = n584_o;
    endcase
  /* project.vhdl:228:48  */
  assign n611_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n611_o)
      2'b00: n612_o = n585_o;
      2'b01: n612_o = n586_o;
      2'b10: n612_o = n587_o;
      2'b11: n612_o = n588_o;
    endcase
  /* project.vhdl:228:48  */
  assign n613_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n613_o)
      2'b00: n614_o = n589_o;
      2'b01: n614_o = n590_o;
      2'b10: n614_o = n591_o;
      2'b11: n614_o = n592_o;
    endcase
  /* project.vhdl:228:48  */
  assign n615_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n615_o)
      2'b00: n616_o = n593_o;
      2'b01: n616_o = n594_o;
      2'b10: n616_o = n595_o;
      2'b11: n616_o = n596_o;
    endcase
  /* project.vhdl:228:48  */
  assign n617_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n617_o)
      2'b00: n618_o = n597_o;
      2'b01: n618_o = n598_o;
      2'b10: n618_o = n599_o;
      2'b11: n618_o = n600_o;
    endcase
  /* project.vhdl:228:48  */
  assign n619_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n619_o)
      2'b00: n620_o = n601_o;
      2'b01: n620_o = n602_o;
      2'b10: n620_o = n603_o;
      2'b11: n620_o = n604_o;
    endcase
  /* project.vhdl:228:48  */
  assign n621_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n621_o)
      2'b00: n622_o = n606_o;
      2'b01: n622_o = n608_o;
      2'b10: n622_o = n610_o;
      2'b11: n622_o = n612_o;
    endcase
  /* project.vhdl:228:48  */
  assign n623_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:228:48  */
  always @*
    case (n623_o)
      2'b00: n624_o = n614_o;
      2'b01: n624_o = n616_o;
      2'b10: n624_o = n618_o;
      2'b11: n624_o = n620_o;
    endcase
  /* project.vhdl:228:48  */
  assign n625_o = i_rom_mrse[4]; // extract
  /* project.vhdl:228:48  */
  assign n626_o = n625_o ? n624_o : n622_o;
  /* project.vhdl:228:48  */
  assign n627_o = rom_mrse[7:0]; // extract
  /* project.vhdl:228:49  */
  assign n628_o = rom_mrse[15:8]; // extract
  assign n629_o = rom_mrse[23:16]; // extract
  assign n630_o = rom_mrse[31:24]; // extract
  assign n631_o = rom_mrse[39:32]; // extract
  assign n632_o = rom_mrse[47:40]; // extract
  assign n633_o = rom_mrse[55:48]; // extract
  assign n634_o = rom_mrse[63:56]; // extract
  assign n635_o = rom_mrse[71:64]; // extract
  assign n636_o = rom_mrse[79:72]; // extract
  assign n637_o = rom_mrse[87:80]; // extract
  assign n638_o = rom_mrse[95:88]; // extract
  assign n639_o = rom_mrse[103:96]; // extract
  assign n640_o = rom_mrse[111:104]; // extract
  assign n641_o = rom_mrse[119:112]; // extract
  assign n642_o = rom_mrse[127:120]; // extract
  assign n643_o = rom_mrse[135:128]; // extract
  assign n644_o = rom_mrse[143:136]; // extract
  assign n645_o = rom_mrse[151:144]; // extract
  assign n646_o = rom_mrse[159:152]; // extract
  assign n647_o = rom_mrse[167:160]; // extract
  assign n648_o = rom_mrse[175:168]; // extract
  assign n649_o = rom_mrse[183:176]; // extract
  assign n650_o = rom_mrse[191:184]; // extract
  assign n651_o = rom_mrse[199:192]; // extract
  assign n652_o = rom_mrse[207:200]; // extract
  assign n653_o = rom_mrse[215:208]; // extract
  assign n654_o = rom_mrse[223:216]; // extract
  assign n655_o = rom_mrse[231:224]; // extract
  assign n656_o = rom_mrse[239:232]; // extract
  assign n657_o = rom_mrse[247:240]; // extract
  assign n658_o = rom_mrse[255:248]; // extract
  /* project.vhdl:246:46  */
  assign n659_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n659_o)
      2'b00: n660_o = n627_o;
      2'b01: n660_o = n628_o;
      2'b10: n660_o = n629_o;
      2'b11: n660_o = n630_o;
    endcase
  /* project.vhdl:246:46  */
  assign n661_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n661_o)
      2'b00: n662_o = n631_o;
      2'b01: n662_o = n632_o;
      2'b10: n662_o = n633_o;
      2'b11: n662_o = n634_o;
    endcase
  /* project.vhdl:246:46  */
  assign n663_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n663_o)
      2'b00: n664_o = n635_o;
      2'b01: n664_o = n636_o;
      2'b10: n664_o = n637_o;
      2'b11: n664_o = n638_o;
    endcase
  /* project.vhdl:246:46  */
  assign n665_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n665_o)
      2'b00: n666_o = n639_o;
      2'b01: n666_o = n640_o;
      2'b10: n666_o = n641_o;
      2'b11: n666_o = n642_o;
    endcase
  /* project.vhdl:246:46  */
  assign n667_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n667_o)
      2'b00: n668_o = n643_o;
      2'b01: n668_o = n644_o;
      2'b10: n668_o = n645_o;
      2'b11: n668_o = n646_o;
    endcase
  /* project.vhdl:246:46  */
  assign n669_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n669_o)
      2'b00: n670_o = n647_o;
      2'b01: n670_o = n648_o;
      2'b10: n670_o = n649_o;
      2'b11: n670_o = n650_o;
    endcase
  /* project.vhdl:246:46  */
  assign n671_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n671_o)
      2'b00: n672_o = n651_o;
      2'b01: n672_o = n652_o;
      2'b10: n672_o = n653_o;
      2'b11: n672_o = n654_o;
    endcase
  /* project.vhdl:246:46  */
  assign n673_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n673_o)
      2'b00: n674_o = n655_o;
      2'b01: n674_o = n656_o;
      2'b10: n674_o = n657_o;
      2'b11: n674_o = n658_o;
    endcase
  /* project.vhdl:246:46  */
  assign n675_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n675_o)
      2'b00: n676_o = n660_o;
      2'b01: n676_o = n662_o;
      2'b10: n676_o = n664_o;
      2'b11: n676_o = n666_o;
    endcase
  /* project.vhdl:246:46  */
  assign n677_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:246:46  */
  always @*
    case (n677_o)
      2'b00: n678_o = n668_o;
      2'b01: n678_o = n670_o;
      2'b10: n678_o = n672_o;
      2'b11: n678_o = n674_o;
    endcase
  /* project.vhdl:246:46  */
  assign n679_o = i_rom_mrse[4]; // extract
  /* project.vhdl:246:46  */
  assign n680_o = n679_o ? n678_o : n676_o;
  /* project.vhdl:247:29  */
  assign n681_o = i_rom_mrse[4]; // extract
  /* project.vhdl:247:29  */
  assign n682_o = ~n681_o;
  /* project.vhdl:247:29  */
  assign n683_o = i_rom_mrse[3]; // extract
  /* project.vhdl:247:29  */
  assign n684_o = ~n683_o;
  /* project.vhdl:247:29  */
  assign n685_o = n682_o & n684_o;
  /* project.vhdl:247:29  */
  assign n686_o = n682_o & n683_o;
  /* project.vhdl:247:29  */
  assign n687_o = n681_o & n684_o;
  /* project.vhdl:247:29  */
  assign n688_o = n681_o & n683_o;
  /* project.vhdl:247:29  */
  assign n689_o = i_rom_mrse[2]; // extract
  /* project.vhdl:247:29  */
  assign n690_o = ~n689_o;
  /* project.vhdl:247:29  */
  assign n691_o = n685_o & n690_o;
  /* project.vhdl:247:29  */
  assign n692_o = n685_o & n689_o;
  /* project.vhdl:247:29  */
  assign n693_o = n686_o & n690_o;
  /* project.vhdl:247:29  */
  assign n694_o = n686_o & n689_o;
  /* project.vhdl:247:29  */
  assign n695_o = n687_o & n690_o;
  /* project.vhdl:247:29  */
  assign n696_o = n687_o & n689_o;
  /* project.vhdl:247:29  */
  assign n697_o = n688_o & n690_o;
  /* project.vhdl:247:29  */
  assign n698_o = n688_o & n689_o;
  /* project.vhdl:247:29  */
  assign n699_o = i_rom_mrse[1]; // extract
  /* project.vhdl:247:29  */
  assign n700_o = ~n699_o;
  /* project.vhdl:247:29  */
  assign n701_o = n691_o & n700_o;
  /* project.vhdl:247:29  */
  assign n702_o = n691_o & n699_o;
  /* project.vhdl:247:29  */
  assign n703_o = n692_o & n700_o;
  /* project.vhdl:247:29  */
  assign n704_o = n692_o & n699_o;
  /* project.vhdl:247:29  */
  assign n705_o = n693_o & n700_o;
  /* project.vhdl:247:29  */
  assign n706_o = n693_o & n699_o;
  /* project.vhdl:247:29  */
  assign n707_o = n694_o & n700_o;
  /* project.vhdl:247:29  */
  assign n708_o = n694_o & n699_o;
  /* project.vhdl:247:29  */
  assign n709_o = n695_o & n700_o;
  /* project.vhdl:247:29  */
  assign n710_o = n695_o & n699_o;
  /* project.vhdl:247:29  */
  assign n711_o = n696_o & n700_o;
  /* project.vhdl:247:29  */
  assign n712_o = n696_o & n699_o;
  /* project.vhdl:247:29  */
  assign n713_o = n697_o & n700_o;
  /* project.vhdl:247:29  */
  assign n714_o = n697_o & n699_o;
  /* project.vhdl:247:29  */
  assign n715_o = n698_o & n700_o;
  /* project.vhdl:247:29  */
  assign n716_o = n698_o & n699_o;
  /* project.vhdl:247:29  */
  assign n717_o = i_rom_mrse[0]; // extract
  /* project.vhdl:247:29  */
  assign n718_o = ~n717_o;
  /* project.vhdl:247:29  */
  assign n719_o = n701_o & n718_o;
  /* project.vhdl:247:29  */
  assign n720_o = n701_o & n717_o;
  /* project.vhdl:247:29  */
  assign n721_o = n702_o & n718_o;
  /* project.vhdl:247:29  */
  assign n722_o = n702_o & n717_o;
  /* project.vhdl:247:29  */
  assign n723_o = n703_o & n718_o;
  /* project.vhdl:247:29  */
  assign n724_o = n703_o & n717_o;
  /* project.vhdl:247:29  */
  assign n725_o = n704_o & n718_o;
  /* project.vhdl:247:29  */
  assign n726_o = n704_o & n717_o;
  /* project.vhdl:247:29  */
  assign n727_o = n705_o & n718_o;
  /* project.vhdl:247:29  */
  assign n728_o = n705_o & n717_o;
  /* project.vhdl:247:29  */
  assign n729_o = n706_o & n718_o;
  /* project.vhdl:247:29  */
  assign n730_o = n706_o & n717_o;
  /* project.vhdl:247:29  */
  assign n731_o = n707_o & n718_o;
  /* project.vhdl:247:29  */
  assign n732_o = n707_o & n717_o;
  /* project.vhdl:247:29  */
  assign n733_o = n708_o & n718_o;
  /* project.vhdl:247:29  */
  assign n734_o = n708_o & n717_o;
  /* project.vhdl:247:29  */
  assign n735_o = n709_o & n718_o;
  /* project.vhdl:247:29  */
  assign n736_o = n709_o & n717_o;
  /* project.vhdl:247:29  */
  assign n737_o = n710_o & n718_o;
  /* project.vhdl:247:29  */
  assign n738_o = n710_o & n717_o;
  /* project.vhdl:247:29  */
  assign n739_o = n711_o & n718_o;
  /* project.vhdl:247:29  */
  assign n740_o = n711_o & n717_o;
  /* project.vhdl:247:29  */
  assign n741_o = n712_o & n718_o;
  /* project.vhdl:247:29  */
  assign n742_o = n712_o & n717_o;
  /* project.vhdl:247:29  */
  assign n743_o = n713_o & n718_o;
  /* project.vhdl:247:29  */
  assign n744_o = n713_o & n717_o;
  /* project.vhdl:247:29  */
  assign n745_o = n714_o & n718_o;
  /* project.vhdl:247:29  */
  assign n746_o = n714_o & n717_o;
  /* project.vhdl:247:29  */
  assign n747_o = n715_o & n718_o;
  /* project.vhdl:247:29  */
  assign n748_o = n715_o & n717_o;
  /* project.vhdl:247:29  */
  assign n749_o = n716_o & n718_o;
  /* project.vhdl:247:29  */
  assign n750_o = n716_o & n717_o;
  assign n751_o = n57_o[7:0]; // extract
  /* project.vhdl:247:29  */
  assign n752_o = n719_o ? n202_o : n751_o;
  assign n753_o = n57_o[15:8]; // extract
  /* project.vhdl:247:29  */
  assign n754_o = n720_o ? n202_o : n753_o;
  assign n755_o = n57_o[23:16]; // extract
  /* project.vhdl:247:29  */
  assign n756_o = n721_o ? n202_o : n755_o;
  assign n757_o = n57_o[31:24]; // extract
  /* project.vhdl:247:29  */
  assign n758_o = n722_o ? n202_o : n757_o;
  assign n759_o = n57_o[39:32]; // extract
  /* project.vhdl:247:29  */
  assign n760_o = n723_o ? n202_o : n759_o;
  assign n761_o = n57_o[47:40]; // extract
  /* project.vhdl:247:29  */
  assign n762_o = n724_o ? n202_o : n761_o;
  assign n763_o = n57_o[55:48]; // extract
  /* project.vhdl:247:29  */
  assign n764_o = n725_o ? n202_o : n763_o;
  assign n765_o = n57_o[63:56]; // extract
  /* project.vhdl:247:29  */
  assign n766_o = n726_o ? n202_o : n765_o;
  assign n767_o = n57_o[71:64]; // extract
  /* project.vhdl:247:29  */
  assign n768_o = n727_o ? n202_o : n767_o;
  assign n769_o = n57_o[79:72]; // extract
  /* project.vhdl:247:29  */
  assign n770_o = n728_o ? n202_o : n769_o;
  assign n771_o = n57_o[87:80]; // extract
  /* project.vhdl:247:29  */
  assign n772_o = n729_o ? n202_o : n771_o;
  assign n773_o = n57_o[95:88]; // extract
  /* project.vhdl:247:29  */
  assign n774_o = n730_o ? n202_o : n773_o;
  assign n775_o = n57_o[103:96]; // extract
  /* project.vhdl:247:29  */
  assign n776_o = n731_o ? n202_o : n775_o;
  assign n777_o = n57_o[111:104]; // extract
  /* project.vhdl:247:29  */
  assign n778_o = n732_o ? n202_o : n777_o;
  assign n779_o = n57_o[119:112]; // extract
  /* project.vhdl:247:29  */
  assign n780_o = n733_o ? n202_o : n779_o;
  assign n781_o = n57_o[127:120]; // extract
  /* project.vhdl:247:29  */
  assign n782_o = n734_o ? n202_o : n781_o;
  assign n783_o = n57_o[135:128]; // extract
  /* project.vhdl:247:29  */
  assign n784_o = n735_o ? n202_o : n783_o;
  assign n785_o = n57_o[143:136]; // extract
  /* project.vhdl:247:29  */
  assign n786_o = n736_o ? n202_o : n785_o;
  assign n787_o = n57_o[151:144]; // extract
  /* project.vhdl:247:29  */
  assign n788_o = n737_o ? n202_o : n787_o;
  assign n789_o = n57_o[159:152]; // extract
  /* project.vhdl:247:29  */
  assign n790_o = n738_o ? n202_o : n789_o;
  assign n791_o = n57_o[167:160]; // extract
  /* project.vhdl:247:29  */
  assign n792_o = n739_o ? n202_o : n791_o;
  assign n793_o = n57_o[175:168]; // extract
  /* project.vhdl:247:29  */
  assign n794_o = n740_o ? n202_o : n793_o;
  assign n795_o = n57_o[183:176]; // extract
  /* project.vhdl:247:29  */
  assign n796_o = n741_o ? n202_o : n795_o;
  assign n797_o = n57_o[191:184]; // extract
  /* project.vhdl:247:29  */
  assign n798_o = n742_o ? n202_o : n797_o;
  assign n799_o = n57_o[199:192]; // extract
  /* project.vhdl:247:29  */
  assign n800_o = n743_o ? n202_o : n799_o;
  assign n801_o = n57_o[207:200]; // extract
  /* project.vhdl:247:29  */
  assign n802_o = n744_o ? n202_o : n801_o;
  assign n803_o = n57_o[215:208]; // extract
  /* project.vhdl:247:29  */
  assign n804_o = n745_o ? n202_o : n803_o;
  assign n805_o = n57_o[223:216]; // extract
  /* project.vhdl:247:29  */
  assign n806_o = n746_o ? n202_o : n805_o;
  assign n807_o = n57_o[231:224]; // extract
  /* project.vhdl:247:29  */
  assign n808_o = n747_o ? n202_o : n807_o;
  assign n809_o = n57_o[239:232]; // extract
  /* project.vhdl:247:29  */
  assign n810_o = n748_o ? n202_o : n809_o;
  assign n811_o = n57_o[247:240]; // extract
  /* project.vhdl:247:29  */
  assign n812_o = n749_o ? n202_o : n811_o;
  assign n813_o = n57_o[255:248]; // extract
  /* project.vhdl:247:29  */
  assign n814_o = n750_o ? n202_o : n813_o;
  assign n815_o = {n814_o, n812_o, n810_o, n808_o, n806_o, n804_o, n802_o, n800_o, n798_o, n796_o, n794_o, n792_o, n790_o, n788_o, n786_o, n784_o, n782_o, n780_o, n778_o, n776_o, n774_o, n772_o, n770_o, n768_o, n766_o, n764_o, n762_o, n760_o, n758_o, n756_o, n754_o, n752_o};
  /* project.vhdl:247:38  */
  assign n816_o = rom_mrse[7:0]; // extract
  /* project.vhdl:247:29  */
  assign n817_o = rom_mrse[15:8]; // extract
  assign n818_o = rom_mrse[23:16]; // extract
  assign n819_o = rom_mrse[31:24]; // extract
  assign n820_o = rom_mrse[39:32]; // extract
  assign n821_o = rom_mrse[47:40]; // extract
  assign n822_o = rom_mrse[55:48]; // extract
  assign n823_o = rom_mrse[63:56]; // extract
  assign n824_o = rom_mrse[71:64]; // extract
  assign n825_o = rom_mrse[79:72]; // extract
  assign n826_o = rom_mrse[87:80]; // extract
  assign n827_o = rom_mrse[95:88]; // extract
  assign n828_o = rom_mrse[103:96]; // extract
  assign n829_o = rom_mrse[111:104]; // extract
  assign n830_o = rom_mrse[119:112]; // extract
  assign n831_o = rom_mrse[127:120]; // extract
  assign n832_o = rom_mrse[135:128]; // extract
  assign n833_o = rom_mrse[143:136]; // extract
  assign n834_o = rom_mrse[151:144]; // extract
  assign n835_o = rom_mrse[159:152]; // extract
  assign n836_o = rom_mrse[167:160]; // extract
  assign n837_o = rom_mrse[175:168]; // extract
  assign n838_o = rom_mrse[183:176]; // extract
  assign n839_o = rom_mrse[191:184]; // extract
  assign n840_o = rom_mrse[199:192]; // extract
  assign n841_o = rom_mrse[207:200]; // extract
  assign n842_o = rom_mrse[215:208]; // extract
  assign n843_o = rom_mrse[223:216]; // extract
  assign n844_o = rom_mrse[231:224]; // extract
  assign n845_o = rom_mrse[239:232]; // extract
  assign n846_o = rom_mrse[247:240]; // extract
  assign n847_o = rom_mrse[255:248]; // extract
  /* project.vhdl:250:48  */
  assign n848_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n848_o)
      2'b00: n849_o = n816_o;
      2'b01: n849_o = n817_o;
      2'b10: n849_o = n818_o;
      2'b11: n849_o = n819_o;
    endcase
  /* project.vhdl:250:48  */
  assign n850_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n850_o)
      2'b00: n851_o = n820_o;
      2'b01: n851_o = n821_o;
      2'b10: n851_o = n822_o;
      2'b11: n851_o = n823_o;
    endcase
  /* project.vhdl:250:48  */
  assign n852_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n852_o)
      2'b00: n853_o = n824_o;
      2'b01: n853_o = n825_o;
      2'b10: n853_o = n826_o;
      2'b11: n853_o = n827_o;
    endcase
  /* project.vhdl:250:48  */
  assign n854_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n854_o)
      2'b00: n855_o = n828_o;
      2'b01: n855_o = n829_o;
      2'b10: n855_o = n830_o;
      2'b11: n855_o = n831_o;
    endcase
  /* project.vhdl:250:48  */
  assign n856_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n856_o)
      2'b00: n857_o = n832_o;
      2'b01: n857_o = n833_o;
      2'b10: n857_o = n834_o;
      2'b11: n857_o = n835_o;
    endcase
  /* project.vhdl:250:48  */
  assign n858_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n858_o)
      2'b00: n859_o = n836_o;
      2'b01: n859_o = n837_o;
      2'b10: n859_o = n838_o;
      2'b11: n859_o = n839_o;
    endcase
  /* project.vhdl:250:48  */
  assign n860_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n860_o)
      2'b00: n861_o = n840_o;
      2'b01: n861_o = n841_o;
      2'b10: n861_o = n842_o;
      2'b11: n861_o = n843_o;
    endcase
  /* project.vhdl:250:48  */
  assign n862_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n862_o)
      2'b00: n863_o = n844_o;
      2'b01: n863_o = n845_o;
      2'b10: n863_o = n846_o;
      2'b11: n863_o = n847_o;
    endcase
  /* project.vhdl:250:48  */
  assign n864_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n864_o)
      2'b00: n865_o = n849_o;
      2'b01: n865_o = n851_o;
      2'b10: n865_o = n853_o;
      2'b11: n865_o = n855_o;
    endcase
  /* project.vhdl:250:48  */
  assign n866_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:250:48  */
  always @*
    case (n866_o)
      2'b00: n867_o = n857_o;
      2'b01: n867_o = n859_o;
      2'b10: n867_o = n861_o;
      2'b11: n867_o = n863_o;
    endcase
  /* project.vhdl:250:48  */
  assign n868_o = i_rom_mrse[4]; // extract
  /* project.vhdl:250:48  */
  assign n869_o = n868_o ? n867_o : n865_o;
  /* project.vhdl:250:48  */
  assign n870_o = rom_mrse[7:0]; // extract
  /* project.vhdl:250:49  */
  assign n871_o = rom_mrse[15:8]; // extract
  assign n872_o = rom_mrse[23:16]; // extract
  assign n873_o = rom_mrse[31:24]; // extract
  assign n874_o = rom_mrse[39:32]; // extract
  assign n875_o = rom_mrse[47:40]; // extract
  assign n876_o = rom_mrse[55:48]; // extract
  assign n877_o = rom_mrse[63:56]; // extract
  assign n878_o = rom_mrse[71:64]; // extract
  assign n879_o = rom_mrse[79:72]; // extract
  assign n880_o = rom_mrse[87:80]; // extract
  assign n881_o = rom_mrse[95:88]; // extract
  assign n882_o = rom_mrse[103:96]; // extract
  assign n883_o = rom_mrse[111:104]; // extract
  assign n884_o = rom_mrse[119:112]; // extract
  assign n885_o = rom_mrse[127:120]; // extract
  assign n886_o = rom_mrse[135:128]; // extract
  assign n887_o = rom_mrse[143:136]; // extract
  assign n888_o = rom_mrse[151:144]; // extract
  assign n889_o = rom_mrse[159:152]; // extract
  assign n890_o = rom_mrse[167:160]; // extract
  assign n891_o = rom_mrse[175:168]; // extract
  assign n892_o = rom_mrse[183:176]; // extract
  assign n893_o = rom_mrse[191:184]; // extract
  assign n894_o = rom_mrse[199:192]; // extract
  assign n895_o = rom_mrse[207:200]; // extract
  assign n896_o = rom_mrse[215:208]; // extract
  assign n897_o = rom_mrse[223:216]; // extract
  assign n898_o = rom_mrse[231:224]; // extract
  assign n899_o = rom_mrse[239:232]; // extract
  assign n900_o = rom_mrse[247:240]; // extract
  assign n901_o = rom_mrse[255:248]; // extract
  /* project.vhdl:259:46  */
  assign n902_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n902_o)
      2'b00: n903_o = n870_o;
      2'b01: n903_o = n871_o;
      2'b10: n903_o = n872_o;
      2'b11: n903_o = n873_o;
    endcase
  /* project.vhdl:259:46  */
  assign n904_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n904_o)
      2'b00: n905_o = n874_o;
      2'b01: n905_o = n875_o;
      2'b10: n905_o = n876_o;
      2'b11: n905_o = n877_o;
    endcase
  /* project.vhdl:259:46  */
  assign n906_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n906_o)
      2'b00: n907_o = n878_o;
      2'b01: n907_o = n879_o;
      2'b10: n907_o = n880_o;
      2'b11: n907_o = n881_o;
    endcase
  /* project.vhdl:259:46  */
  assign n908_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n908_o)
      2'b00: n909_o = n882_o;
      2'b01: n909_o = n883_o;
      2'b10: n909_o = n884_o;
      2'b11: n909_o = n885_o;
    endcase
  /* project.vhdl:259:46  */
  assign n910_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n910_o)
      2'b00: n911_o = n886_o;
      2'b01: n911_o = n887_o;
      2'b10: n911_o = n888_o;
      2'b11: n911_o = n889_o;
    endcase
  /* project.vhdl:259:46  */
  assign n912_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n912_o)
      2'b00: n913_o = n890_o;
      2'b01: n913_o = n891_o;
      2'b10: n913_o = n892_o;
      2'b11: n913_o = n893_o;
    endcase
  /* project.vhdl:259:46  */
  assign n914_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n914_o)
      2'b00: n915_o = n894_o;
      2'b01: n915_o = n895_o;
      2'b10: n915_o = n896_o;
      2'b11: n915_o = n897_o;
    endcase
  /* project.vhdl:259:46  */
  assign n916_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n916_o)
      2'b00: n917_o = n898_o;
      2'b01: n917_o = n899_o;
      2'b10: n917_o = n900_o;
      2'b11: n917_o = n901_o;
    endcase
  /* project.vhdl:259:46  */
  assign n918_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n918_o)
      2'b00: n919_o = n903_o;
      2'b01: n919_o = n905_o;
      2'b10: n919_o = n907_o;
      2'b11: n919_o = n909_o;
    endcase
  /* project.vhdl:259:46  */
  assign n920_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:259:46  */
  always @*
    case (n920_o)
      2'b00: n921_o = n911_o;
      2'b01: n921_o = n913_o;
      2'b10: n921_o = n915_o;
      2'b11: n921_o = n917_o;
    endcase
  /* project.vhdl:259:46  */
  assign n922_o = i_rom_mrse[4]; // extract
  /* project.vhdl:259:46  */
  assign n923_o = n922_o ? n921_o : n919_o;
  /* project.vhdl:260:29  */
  assign n924_o = i_rom_mrse[4]; // extract
  /* project.vhdl:260:29  */
  assign n925_o = ~n924_o;
  /* project.vhdl:260:29  */
  assign n926_o = i_rom_mrse[3]; // extract
  /* project.vhdl:260:29  */
  assign n927_o = ~n926_o;
  /* project.vhdl:260:29  */
  assign n928_o = n925_o & n927_o;
  /* project.vhdl:260:29  */
  assign n929_o = n925_o & n926_o;
  /* project.vhdl:260:29  */
  assign n930_o = n924_o & n927_o;
  /* project.vhdl:260:29  */
  assign n931_o = n924_o & n926_o;
  /* project.vhdl:260:29  */
  assign n932_o = i_rom_mrse[2]; // extract
  /* project.vhdl:260:29  */
  assign n933_o = ~n932_o;
  /* project.vhdl:260:29  */
  assign n934_o = n928_o & n933_o;
  /* project.vhdl:260:29  */
  assign n935_o = n928_o & n932_o;
  /* project.vhdl:260:29  */
  assign n936_o = n929_o & n933_o;
  /* project.vhdl:260:29  */
  assign n937_o = n929_o & n932_o;
  /* project.vhdl:260:29  */
  assign n938_o = n930_o & n933_o;
  /* project.vhdl:260:29  */
  assign n939_o = n930_o & n932_o;
  /* project.vhdl:260:29  */
  assign n940_o = n931_o & n933_o;
  /* project.vhdl:260:29  */
  assign n941_o = n931_o & n932_o;
  /* project.vhdl:260:29  */
  assign n942_o = i_rom_mrse[1]; // extract
  /* project.vhdl:260:29  */
  assign n943_o = ~n942_o;
  /* project.vhdl:260:29  */
  assign n944_o = n934_o & n943_o;
  /* project.vhdl:260:29  */
  assign n945_o = n934_o & n942_o;
  /* project.vhdl:260:29  */
  assign n946_o = n935_o & n943_o;
  /* project.vhdl:260:29  */
  assign n947_o = n935_o & n942_o;
  /* project.vhdl:260:29  */
  assign n948_o = n936_o & n943_o;
  /* project.vhdl:260:29  */
  assign n949_o = n936_o & n942_o;
  /* project.vhdl:260:29  */
  assign n950_o = n937_o & n943_o;
  /* project.vhdl:260:29  */
  assign n951_o = n937_o & n942_o;
  /* project.vhdl:260:29  */
  assign n952_o = n938_o & n943_o;
  /* project.vhdl:260:29  */
  assign n953_o = n938_o & n942_o;
  /* project.vhdl:260:29  */
  assign n954_o = n939_o & n943_o;
  /* project.vhdl:260:29  */
  assign n955_o = n939_o & n942_o;
  /* project.vhdl:260:29  */
  assign n956_o = n940_o & n943_o;
  /* project.vhdl:260:29  */
  assign n957_o = n940_o & n942_o;
  /* project.vhdl:260:29  */
  assign n958_o = n941_o & n943_o;
  /* project.vhdl:260:29  */
  assign n959_o = n941_o & n942_o;
  /* project.vhdl:260:29  */
  assign n960_o = i_rom_mrse[0]; // extract
  /* project.vhdl:260:29  */
  assign n961_o = ~n960_o;
  /* project.vhdl:260:29  */
  assign n962_o = n944_o & n961_o;
  /* project.vhdl:260:29  */
  assign n963_o = n944_o & n960_o;
  /* project.vhdl:260:29  */
  assign n964_o = n945_o & n961_o;
  /* project.vhdl:260:29  */
  assign n965_o = n945_o & n960_o;
  /* project.vhdl:260:29  */
  assign n966_o = n946_o & n961_o;
  /* project.vhdl:260:29  */
  assign n967_o = n946_o & n960_o;
  /* project.vhdl:260:29  */
  assign n968_o = n947_o & n961_o;
  /* project.vhdl:260:29  */
  assign n969_o = n947_o & n960_o;
  /* project.vhdl:260:29  */
  assign n970_o = n948_o & n961_o;
  /* project.vhdl:260:29  */
  assign n971_o = n948_o & n960_o;
  /* project.vhdl:260:29  */
  assign n972_o = n949_o & n961_o;
  /* project.vhdl:260:29  */
  assign n973_o = n949_o & n960_o;
  /* project.vhdl:260:29  */
  assign n974_o = n950_o & n961_o;
  /* project.vhdl:260:29  */
  assign n975_o = n950_o & n960_o;
  /* project.vhdl:260:29  */
  assign n976_o = n951_o & n961_o;
  /* project.vhdl:260:29  */
  assign n977_o = n951_o & n960_o;
  /* project.vhdl:260:29  */
  assign n978_o = n952_o & n961_o;
  /* project.vhdl:260:29  */
  assign n979_o = n952_o & n960_o;
  /* project.vhdl:260:29  */
  assign n980_o = n953_o & n961_o;
  /* project.vhdl:260:29  */
  assign n981_o = n953_o & n960_o;
  /* project.vhdl:260:29  */
  assign n982_o = n954_o & n961_o;
  /* project.vhdl:260:29  */
  assign n983_o = n954_o & n960_o;
  /* project.vhdl:260:29  */
  assign n984_o = n955_o & n961_o;
  /* project.vhdl:260:29  */
  assign n985_o = n955_o & n960_o;
  /* project.vhdl:260:29  */
  assign n986_o = n956_o & n961_o;
  /* project.vhdl:260:29  */
  assign n987_o = n956_o & n960_o;
  /* project.vhdl:260:29  */
  assign n988_o = n957_o & n961_o;
  /* project.vhdl:260:29  */
  assign n989_o = n957_o & n960_o;
  /* project.vhdl:260:29  */
  assign n990_o = n958_o & n961_o;
  /* project.vhdl:260:29  */
  assign n991_o = n958_o & n960_o;
  /* project.vhdl:260:29  */
  assign n992_o = n959_o & n961_o;
  /* project.vhdl:260:29  */
  assign n993_o = n959_o & n960_o;
  assign n994_o = n57_o[7:0]; // extract
  /* project.vhdl:260:29  */
  assign n995_o = n962_o ? n228_o : n994_o;
  assign n996_o = n57_o[15:8]; // extract
  /* project.vhdl:260:29  */
  assign n997_o = n963_o ? n228_o : n996_o;
  assign n998_o = n57_o[23:16]; // extract
  /* project.vhdl:260:29  */
  assign n999_o = n964_o ? n228_o : n998_o;
  assign n1000_o = n57_o[31:24]; // extract
  /* project.vhdl:260:29  */
  assign n1001_o = n965_o ? n228_o : n1000_o;
  assign n1002_o = n57_o[39:32]; // extract
  /* project.vhdl:260:29  */
  assign n1003_o = n966_o ? n228_o : n1002_o;
  assign n1004_o = n57_o[47:40]; // extract
  /* project.vhdl:260:29  */
  assign n1005_o = n967_o ? n228_o : n1004_o;
  assign n1006_o = n57_o[55:48]; // extract
  /* project.vhdl:260:29  */
  assign n1007_o = n968_o ? n228_o : n1006_o;
  assign n1008_o = n57_o[63:56]; // extract
  /* project.vhdl:260:29  */
  assign n1009_o = n969_o ? n228_o : n1008_o;
  assign n1010_o = n57_o[71:64]; // extract
  /* project.vhdl:260:29  */
  assign n1011_o = n970_o ? n228_o : n1010_o;
  assign n1012_o = n57_o[79:72]; // extract
  /* project.vhdl:260:29  */
  assign n1013_o = n971_o ? n228_o : n1012_o;
  assign n1014_o = n57_o[87:80]; // extract
  /* project.vhdl:260:29  */
  assign n1015_o = n972_o ? n228_o : n1014_o;
  assign n1016_o = n57_o[95:88]; // extract
  /* project.vhdl:260:29  */
  assign n1017_o = n973_o ? n228_o : n1016_o;
  assign n1018_o = n57_o[103:96]; // extract
  /* project.vhdl:260:29  */
  assign n1019_o = n974_o ? n228_o : n1018_o;
  assign n1020_o = n57_o[111:104]; // extract
  /* project.vhdl:260:29  */
  assign n1021_o = n975_o ? n228_o : n1020_o;
  assign n1022_o = n57_o[119:112]; // extract
  /* project.vhdl:260:29  */
  assign n1023_o = n976_o ? n228_o : n1022_o;
  assign n1024_o = n57_o[127:120]; // extract
  /* project.vhdl:260:29  */
  assign n1025_o = n977_o ? n228_o : n1024_o;
  assign n1026_o = n57_o[135:128]; // extract
  /* project.vhdl:260:29  */
  assign n1027_o = n978_o ? n228_o : n1026_o;
  assign n1028_o = n57_o[143:136]; // extract
  /* project.vhdl:260:29  */
  assign n1029_o = n979_o ? n228_o : n1028_o;
  assign n1030_o = n57_o[151:144]; // extract
  /* project.vhdl:260:29  */
  assign n1031_o = n980_o ? n228_o : n1030_o;
  assign n1032_o = n57_o[159:152]; // extract
  /* project.vhdl:260:29  */
  assign n1033_o = n981_o ? n228_o : n1032_o;
  assign n1034_o = n57_o[167:160]; // extract
  /* project.vhdl:260:29  */
  assign n1035_o = n982_o ? n228_o : n1034_o;
  assign n1036_o = n57_o[175:168]; // extract
  /* project.vhdl:260:29  */
  assign n1037_o = n983_o ? n228_o : n1036_o;
  assign n1038_o = n57_o[183:176]; // extract
  /* project.vhdl:260:29  */
  assign n1039_o = n984_o ? n228_o : n1038_o;
  assign n1040_o = n57_o[191:184]; // extract
  /* project.vhdl:260:29  */
  assign n1041_o = n985_o ? n228_o : n1040_o;
  assign n1042_o = n57_o[199:192]; // extract
  /* project.vhdl:260:29  */
  assign n1043_o = n986_o ? n228_o : n1042_o;
  assign n1044_o = n57_o[207:200]; // extract
  /* project.vhdl:260:29  */
  assign n1045_o = n987_o ? n228_o : n1044_o;
  assign n1046_o = n57_o[215:208]; // extract
  /* project.vhdl:260:29  */
  assign n1047_o = n988_o ? n228_o : n1046_o;
  assign n1048_o = n57_o[223:216]; // extract
  /* project.vhdl:260:29  */
  assign n1049_o = n989_o ? n228_o : n1048_o;
  assign n1050_o = n57_o[231:224]; // extract
  /* project.vhdl:260:29  */
  assign n1051_o = n990_o ? n228_o : n1050_o;
  assign n1052_o = n57_o[239:232]; // extract
  /* project.vhdl:260:29  */
  assign n1053_o = n991_o ? n228_o : n1052_o;
  assign n1054_o = n57_o[247:240]; // extract
  /* project.vhdl:260:29  */
  assign n1055_o = n992_o ? n228_o : n1054_o;
  assign n1056_o = n57_o[255:248]; // extract
  /* project.vhdl:260:29  */
  assign n1057_o = n993_o ? n228_o : n1056_o;
  assign n1058_o = {n1057_o, n1055_o, n1053_o, n1051_o, n1049_o, n1047_o, n1045_o, n1043_o, n1041_o, n1039_o, n1037_o, n1035_o, n1033_o, n1031_o, n1029_o, n1027_o, n1025_o, n1023_o, n1021_o, n1019_o, n1017_o, n1015_o, n1013_o, n1011_o, n1009_o, n1007_o, n1005_o, n1003_o, n1001_o, n999_o, n997_o, n995_o};
  /* project.vhdl:260:38  */
  assign n1059_o = rom_mrse[7:0]; // extract
  /* project.vhdl:260:29  */
  assign n1060_o = rom_mrse[15:8]; // extract
  assign n1061_o = rom_mrse[23:16]; // extract
  assign n1062_o = rom_mrse[31:24]; // extract
  assign n1063_o = rom_mrse[39:32]; // extract
  assign n1064_o = rom_mrse[47:40]; // extract
  assign n1065_o = rom_mrse[55:48]; // extract
  assign n1066_o = rom_mrse[63:56]; // extract
  assign n1067_o = rom_mrse[71:64]; // extract
  assign n1068_o = rom_mrse[79:72]; // extract
  assign n1069_o = rom_mrse[87:80]; // extract
  assign n1070_o = rom_mrse[95:88]; // extract
  assign n1071_o = rom_mrse[103:96]; // extract
  assign n1072_o = rom_mrse[111:104]; // extract
  assign n1073_o = rom_mrse[119:112]; // extract
  assign n1074_o = rom_mrse[127:120]; // extract
  assign n1075_o = rom_mrse[135:128]; // extract
  assign n1076_o = rom_mrse[143:136]; // extract
  assign n1077_o = rom_mrse[151:144]; // extract
  assign n1078_o = rom_mrse[159:152]; // extract
  assign n1079_o = rom_mrse[167:160]; // extract
  assign n1080_o = rom_mrse[175:168]; // extract
  assign n1081_o = rom_mrse[183:176]; // extract
  assign n1082_o = rom_mrse[191:184]; // extract
  assign n1083_o = rom_mrse[199:192]; // extract
  assign n1084_o = rom_mrse[207:200]; // extract
  assign n1085_o = rom_mrse[215:208]; // extract
  assign n1086_o = rom_mrse[223:216]; // extract
  assign n1087_o = rom_mrse[231:224]; // extract
  assign n1088_o = rom_mrse[239:232]; // extract
  assign n1089_o = rom_mrse[247:240]; // extract
  assign n1090_o = rom_mrse[255:248]; // extract
  /* project.vhdl:263:48  */
  assign n1091_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1091_o)
      2'b00: n1092_o = n1059_o;
      2'b01: n1092_o = n1060_o;
      2'b10: n1092_o = n1061_o;
      2'b11: n1092_o = n1062_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1093_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1093_o)
      2'b00: n1094_o = n1063_o;
      2'b01: n1094_o = n1064_o;
      2'b10: n1094_o = n1065_o;
      2'b11: n1094_o = n1066_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1095_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1095_o)
      2'b00: n1096_o = n1067_o;
      2'b01: n1096_o = n1068_o;
      2'b10: n1096_o = n1069_o;
      2'b11: n1096_o = n1070_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1097_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1097_o)
      2'b00: n1098_o = n1071_o;
      2'b01: n1098_o = n1072_o;
      2'b10: n1098_o = n1073_o;
      2'b11: n1098_o = n1074_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1099_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1099_o)
      2'b00: n1100_o = n1075_o;
      2'b01: n1100_o = n1076_o;
      2'b10: n1100_o = n1077_o;
      2'b11: n1100_o = n1078_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1101_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1101_o)
      2'b00: n1102_o = n1079_o;
      2'b01: n1102_o = n1080_o;
      2'b10: n1102_o = n1081_o;
      2'b11: n1102_o = n1082_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1103_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1103_o)
      2'b00: n1104_o = n1083_o;
      2'b01: n1104_o = n1084_o;
      2'b10: n1104_o = n1085_o;
      2'b11: n1104_o = n1086_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1105_o = i_rom_mrse[1:0]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1105_o)
      2'b00: n1106_o = n1087_o;
      2'b01: n1106_o = n1088_o;
      2'b10: n1106_o = n1089_o;
      2'b11: n1106_o = n1090_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1107_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1107_o)
      2'b00: n1108_o = n1092_o;
      2'b01: n1108_o = n1094_o;
      2'b10: n1108_o = n1096_o;
      2'b11: n1108_o = n1098_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1109_o = i_rom_mrse[3:2]; // extract
  /* project.vhdl:263:48  */
  always @*
    case (n1109_o)
      2'b00: n1110_o = n1100_o;
      2'b01: n1110_o = n1102_o;
      2'b10: n1110_o = n1104_o;
      2'b11: n1110_o = n1106_o;
    endcase
  /* project.vhdl:263:48  */
  assign n1111_o = i_rom_mrse[4]; // extract
  /* project.vhdl:263:48  */
  assign n1112_o = n1111_o ? n1110_o : n1108_o;
endmodule

